module tt_um_ashleyjr_delay_line (VGND,
    VPWR,
    clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input VGND;
 input VPWR;
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire net1;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net2;
 wire net3;
 wire net4;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net5;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net6;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire \u_delay_line.bulk_0 ;
 wire \u_delay_line.bulk_1 ;
 wire \u_delay_line.bulk_10 ;
 wire \u_delay_line.bulk_11 ;
 wire \u_delay_line.bulk_12 ;
 wire \u_delay_line.bulk_13 ;
 wire \u_delay_line.bulk_14 ;
 wire \u_delay_line.bulk_15 ;
 wire \u_delay_line.bulk_16 ;
 wire \u_delay_line.bulk_17 ;
 wire \u_delay_line.bulk_18 ;
 wire \u_delay_line.bulk_19 ;
 wire \u_delay_line.bulk_2 ;
 wire \u_delay_line.bulk_20 ;
 wire \u_delay_line.bulk_3 ;
 wire \u_delay_line.bulk_4 ;
 wire \u_delay_line.bulk_5 ;
 wire \u_delay_line.bulk_6 ;
 wire \u_delay_line.bulk_7 ;
 wire \u_delay_line.bulk_8 ;
 wire \u_delay_line.bulk_9 ;
 wire \u_delay_line.data_0 ;
 wire \u_delay_line.data_1 ;
 wire \u_delay_line.data_10 ;
 wire \u_delay_line.data_11 ;
 wire \u_delay_line.data_12 ;
 wire \u_delay_line.data_13 ;
 wire \u_delay_line.data_14 ;
 wire \u_delay_line.data_15 ;
 wire \u_delay_line.data_16 ;
 wire \u_delay_line.data_17 ;
 wire \u_delay_line.data_18 ;
 wire \u_delay_line.data_19 ;
 wire \u_delay_line.data_2 ;
 wire \u_delay_line.data_20 ;
 wire \u_delay_line.data_21 ;
 wire \u_delay_line.data_22 ;
 wire \u_delay_line.data_23 ;
 wire \u_delay_line.data_24 ;
 wire \u_delay_line.data_25 ;
 wire \u_delay_line.data_26 ;
 wire \u_delay_line.data_27 ;
 wire \u_delay_line.data_28 ;
 wire \u_delay_line.data_29 ;
 wire \u_delay_line.data_3 ;
 wire \u_delay_line.data_30 ;
 wire \u_delay_line.data_31 ;
 wire \u_delay_line.data_4 ;
 wire \u_delay_line.data_5 ;
 wire \u_delay_line.data_6 ;
 wire \u_delay_line.data_7 ;
 wire \u_delay_line.data_8 ;
 wire \u_delay_line.data_9 ;
 wire \u_delay_line.dl_0 ;
 wire \u_delay_line.dl_1 ;
 wire \u_delay_line.dl_10 ;
 wire \u_delay_line.dl_11 ;
 wire \u_delay_line.dl_12 ;
 wire \u_delay_line.dl_13 ;
 wire \u_delay_line.dl_14 ;
 wire \u_delay_line.dl_15 ;
 wire \u_delay_line.dl_16 ;
 wire \u_delay_line.dl_17 ;
 wire \u_delay_line.dl_18 ;
 wire \u_delay_line.dl_19 ;
 wire \u_delay_line.dl_2 ;
 wire \u_delay_line.dl_20 ;
 wire \u_delay_line.dl_21 ;
 wire \u_delay_line.dl_22 ;
 wire \u_delay_line.dl_23 ;
 wire \u_delay_line.dl_24 ;
 wire \u_delay_line.dl_25 ;
 wire \u_delay_line.dl_26 ;
 wire \u_delay_line.dl_27 ;
 wire \u_delay_line.dl_28 ;
 wire \u_delay_line.dl_29 ;
 wire \u_delay_line.dl_3 ;
 wire \u_delay_line.dl_30 ;
 wire \u_delay_line.dl_31 ;
 wire \u_delay_line.dl_32 ;
 wire \u_delay_line.dl_4 ;
 wire \u_delay_line.dl_5 ;
 wire \u_delay_line.dl_6 ;
 wire \u_delay_line.dl_7 ;
 wire \u_delay_line.dl_8 ;
 wire \u_delay_line.dl_9 ;
 wire \u_delay_line.start_d ;
 wire \u_delay_line.start_q ;
 wire \u_delay_line.u_bulk_0.dl_0 ;
 wire \u_delay_line.u_bulk_0.dl_1 ;
 wire \u_delay_line.u_bulk_0.dl_10 ;
 wire \u_delay_line.u_bulk_0.dl_11 ;
 wire \u_delay_line.u_bulk_0.dl_12 ;
 wire \u_delay_line.u_bulk_0.dl_13 ;
 wire \u_delay_line.u_bulk_0.dl_14 ;
 wire \u_delay_line.u_bulk_0.dl_2 ;
 wire \u_delay_line.u_bulk_0.dl_3 ;
 wire \u_delay_line.u_bulk_0.dl_4 ;
 wire \u_delay_line.u_bulk_0.dl_5 ;
 wire \u_delay_line.u_bulk_0.dl_6 ;
 wire \u_delay_line.u_bulk_0.dl_7 ;
 wire \u_delay_line.u_bulk_0.dl_8 ;
 wire \u_delay_line.u_bulk_0.dl_9 ;
 wire \u_delay_line.u_bulk_1.dl_0 ;
 wire \u_delay_line.u_bulk_1.dl_1 ;
 wire \u_delay_line.u_bulk_1.dl_10 ;
 wire \u_delay_line.u_bulk_1.dl_11 ;
 wire \u_delay_line.u_bulk_1.dl_12 ;
 wire \u_delay_line.u_bulk_1.dl_13 ;
 wire \u_delay_line.u_bulk_1.dl_14 ;
 wire \u_delay_line.u_bulk_1.dl_2 ;
 wire \u_delay_line.u_bulk_1.dl_3 ;
 wire \u_delay_line.u_bulk_1.dl_4 ;
 wire \u_delay_line.u_bulk_1.dl_5 ;
 wire \u_delay_line.u_bulk_1.dl_6 ;
 wire \u_delay_line.u_bulk_1.dl_7 ;
 wire \u_delay_line.u_bulk_1.dl_8 ;
 wire \u_delay_line.u_bulk_1.dl_9 ;
 wire \u_delay_line.u_bulk_10.dl_0 ;
 wire \u_delay_line.u_bulk_10.dl_1 ;
 wire \u_delay_line.u_bulk_10.dl_10 ;
 wire \u_delay_line.u_bulk_10.dl_11 ;
 wire \u_delay_line.u_bulk_10.dl_12 ;
 wire \u_delay_line.u_bulk_10.dl_13 ;
 wire \u_delay_line.u_bulk_10.dl_14 ;
 wire \u_delay_line.u_bulk_10.dl_2 ;
 wire \u_delay_line.u_bulk_10.dl_3 ;
 wire \u_delay_line.u_bulk_10.dl_4 ;
 wire \u_delay_line.u_bulk_10.dl_5 ;
 wire \u_delay_line.u_bulk_10.dl_6 ;
 wire \u_delay_line.u_bulk_10.dl_7 ;
 wire \u_delay_line.u_bulk_10.dl_8 ;
 wire \u_delay_line.u_bulk_10.dl_9 ;
 wire \u_delay_line.u_bulk_11.dl_0 ;
 wire \u_delay_line.u_bulk_11.dl_1 ;
 wire \u_delay_line.u_bulk_11.dl_10 ;
 wire \u_delay_line.u_bulk_11.dl_11 ;
 wire \u_delay_line.u_bulk_11.dl_12 ;
 wire \u_delay_line.u_bulk_11.dl_13 ;
 wire \u_delay_line.u_bulk_11.dl_14 ;
 wire \u_delay_line.u_bulk_11.dl_2 ;
 wire \u_delay_line.u_bulk_11.dl_3 ;
 wire \u_delay_line.u_bulk_11.dl_4 ;
 wire \u_delay_line.u_bulk_11.dl_5 ;
 wire \u_delay_line.u_bulk_11.dl_6 ;
 wire \u_delay_line.u_bulk_11.dl_7 ;
 wire \u_delay_line.u_bulk_11.dl_8 ;
 wire \u_delay_line.u_bulk_11.dl_9 ;
 wire \u_delay_line.u_bulk_12.dl_0 ;
 wire \u_delay_line.u_bulk_12.dl_1 ;
 wire \u_delay_line.u_bulk_12.dl_10 ;
 wire \u_delay_line.u_bulk_12.dl_11 ;
 wire \u_delay_line.u_bulk_12.dl_12 ;
 wire \u_delay_line.u_bulk_12.dl_13 ;
 wire \u_delay_line.u_bulk_12.dl_14 ;
 wire \u_delay_line.u_bulk_12.dl_2 ;
 wire \u_delay_line.u_bulk_12.dl_3 ;
 wire \u_delay_line.u_bulk_12.dl_4 ;
 wire \u_delay_line.u_bulk_12.dl_5 ;
 wire \u_delay_line.u_bulk_12.dl_6 ;
 wire \u_delay_line.u_bulk_12.dl_7 ;
 wire \u_delay_line.u_bulk_12.dl_8 ;
 wire \u_delay_line.u_bulk_12.dl_9 ;
 wire \u_delay_line.u_bulk_13.dl_0 ;
 wire \u_delay_line.u_bulk_13.dl_1 ;
 wire \u_delay_line.u_bulk_13.dl_10 ;
 wire \u_delay_line.u_bulk_13.dl_11 ;
 wire \u_delay_line.u_bulk_13.dl_12 ;
 wire \u_delay_line.u_bulk_13.dl_13 ;
 wire \u_delay_line.u_bulk_13.dl_14 ;
 wire \u_delay_line.u_bulk_13.dl_2 ;
 wire \u_delay_line.u_bulk_13.dl_3 ;
 wire \u_delay_line.u_bulk_13.dl_4 ;
 wire \u_delay_line.u_bulk_13.dl_5 ;
 wire \u_delay_line.u_bulk_13.dl_6 ;
 wire \u_delay_line.u_bulk_13.dl_7 ;
 wire \u_delay_line.u_bulk_13.dl_8 ;
 wire \u_delay_line.u_bulk_13.dl_9 ;
 wire \u_delay_line.u_bulk_14.dl_0 ;
 wire \u_delay_line.u_bulk_14.dl_1 ;
 wire \u_delay_line.u_bulk_14.dl_10 ;
 wire \u_delay_line.u_bulk_14.dl_11 ;
 wire \u_delay_line.u_bulk_14.dl_12 ;
 wire \u_delay_line.u_bulk_14.dl_13 ;
 wire \u_delay_line.u_bulk_14.dl_14 ;
 wire \u_delay_line.u_bulk_14.dl_2 ;
 wire \u_delay_line.u_bulk_14.dl_3 ;
 wire \u_delay_line.u_bulk_14.dl_4 ;
 wire \u_delay_line.u_bulk_14.dl_5 ;
 wire \u_delay_line.u_bulk_14.dl_6 ;
 wire \u_delay_line.u_bulk_14.dl_7 ;
 wire \u_delay_line.u_bulk_14.dl_8 ;
 wire \u_delay_line.u_bulk_14.dl_9 ;
 wire \u_delay_line.u_bulk_15.dl_0 ;
 wire \u_delay_line.u_bulk_15.dl_1 ;
 wire \u_delay_line.u_bulk_15.dl_10 ;
 wire \u_delay_line.u_bulk_15.dl_11 ;
 wire \u_delay_line.u_bulk_15.dl_12 ;
 wire \u_delay_line.u_bulk_15.dl_13 ;
 wire \u_delay_line.u_bulk_15.dl_14 ;
 wire \u_delay_line.u_bulk_15.dl_2 ;
 wire \u_delay_line.u_bulk_15.dl_3 ;
 wire \u_delay_line.u_bulk_15.dl_4 ;
 wire \u_delay_line.u_bulk_15.dl_5 ;
 wire \u_delay_line.u_bulk_15.dl_6 ;
 wire \u_delay_line.u_bulk_15.dl_7 ;
 wire \u_delay_line.u_bulk_15.dl_8 ;
 wire \u_delay_line.u_bulk_15.dl_9 ;
 wire \u_delay_line.u_bulk_16.dl_0 ;
 wire \u_delay_line.u_bulk_16.dl_1 ;
 wire \u_delay_line.u_bulk_16.dl_10 ;
 wire \u_delay_line.u_bulk_16.dl_11 ;
 wire \u_delay_line.u_bulk_16.dl_12 ;
 wire \u_delay_line.u_bulk_16.dl_13 ;
 wire \u_delay_line.u_bulk_16.dl_14 ;
 wire \u_delay_line.u_bulk_16.dl_2 ;
 wire \u_delay_line.u_bulk_16.dl_3 ;
 wire \u_delay_line.u_bulk_16.dl_4 ;
 wire \u_delay_line.u_bulk_16.dl_5 ;
 wire \u_delay_line.u_bulk_16.dl_6 ;
 wire \u_delay_line.u_bulk_16.dl_7 ;
 wire \u_delay_line.u_bulk_16.dl_8 ;
 wire \u_delay_line.u_bulk_16.dl_9 ;
 wire \u_delay_line.u_bulk_17.dl_0 ;
 wire \u_delay_line.u_bulk_17.dl_1 ;
 wire \u_delay_line.u_bulk_17.dl_10 ;
 wire \u_delay_line.u_bulk_17.dl_11 ;
 wire \u_delay_line.u_bulk_17.dl_12 ;
 wire \u_delay_line.u_bulk_17.dl_13 ;
 wire \u_delay_line.u_bulk_17.dl_14 ;
 wire \u_delay_line.u_bulk_17.dl_2 ;
 wire \u_delay_line.u_bulk_17.dl_3 ;
 wire \u_delay_line.u_bulk_17.dl_4 ;
 wire \u_delay_line.u_bulk_17.dl_5 ;
 wire \u_delay_line.u_bulk_17.dl_6 ;
 wire \u_delay_line.u_bulk_17.dl_7 ;
 wire \u_delay_line.u_bulk_17.dl_8 ;
 wire \u_delay_line.u_bulk_17.dl_9 ;
 wire \u_delay_line.u_bulk_18.dl_0 ;
 wire \u_delay_line.u_bulk_18.dl_1 ;
 wire \u_delay_line.u_bulk_18.dl_10 ;
 wire \u_delay_line.u_bulk_18.dl_11 ;
 wire \u_delay_line.u_bulk_18.dl_12 ;
 wire \u_delay_line.u_bulk_18.dl_13 ;
 wire \u_delay_line.u_bulk_18.dl_14 ;
 wire \u_delay_line.u_bulk_18.dl_2 ;
 wire \u_delay_line.u_bulk_18.dl_3 ;
 wire \u_delay_line.u_bulk_18.dl_4 ;
 wire \u_delay_line.u_bulk_18.dl_5 ;
 wire \u_delay_line.u_bulk_18.dl_6 ;
 wire \u_delay_line.u_bulk_18.dl_7 ;
 wire \u_delay_line.u_bulk_18.dl_8 ;
 wire \u_delay_line.u_bulk_18.dl_9 ;
 wire \u_delay_line.u_bulk_19.dl_0 ;
 wire \u_delay_line.u_bulk_19.dl_1 ;
 wire \u_delay_line.u_bulk_19.dl_10 ;
 wire \u_delay_line.u_bulk_19.dl_11 ;
 wire \u_delay_line.u_bulk_19.dl_12 ;
 wire \u_delay_line.u_bulk_19.dl_13 ;
 wire \u_delay_line.u_bulk_19.dl_14 ;
 wire \u_delay_line.u_bulk_19.dl_2 ;
 wire \u_delay_line.u_bulk_19.dl_3 ;
 wire \u_delay_line.u_bulk_19.dl_4 ;
 wire \u_delay_line.u_bulk_19.dl_5 ;
 wire \u_delay_line.u_bulk_19.dl_6 ;
 wire \u_delay_line.u_bulk_19.dl_7 ;
 wire \u_delay_line.u_bulk_19.dl_8 ;
 wire \u_delay_line.u_bulk_19.dl_9 ;
 wire \u_delay_line.u_bulk_2.dl_0 ;
 wire \u_delay_line.u_bulk_2.dl_1 ;
 wire \u_delay_line.u_bulk_2.dl_10 ;
 wire \u_delay_line.u_bulk_2.dl_11 ;
 wire \u_delay_line.u_bulk_2.dl_12 ;
 wire \u_delay_line.u_bulk_2.dl_13 ;
 wire \u_delay_line.u_bulk_2.dl_14 ;
 wire \u_delay_line.u_bulk_2.dl_2 ;
 wire \u_delay_line.u_bulk_2.dl_3 ;
 wire \u_delay_line.u_bulk_2.dl_4 ;
 wire \u_delay_line.u_bulk_2.dl_5 ;
 wire \u_delay_line.u_bulk_2.dl_6 ;
 wire \u_delay_line.u_bulk_2.dl_7 ;
 wire \u_delay_line.u_bulk_2.dl_8 ;
 wire \u_delay_line.u_bulk_2.dl_9 ;
 wire \u_delay_line.u_bulk_20.dl_0 ;
 wire \u_delay_line.u_bulk_20.dl_1 ;
 wire \u_delay_line.u_bulk_20.dl_10 ;
 wire \u_delay_line.u_bulk_20.dl_11 ;
 wire \u_delay_line.u_bulk_20.dl_12 ;
 wire \u_delay_line.u_bulk_20.dl_13 ;
 wire \u_delay_line.u_bulk_20.dl_14 ;
 wire \u_delay_line.u_bulk_20.dl_2 ;
 wire \u_delay_line.u_bulk_20.dl_3 ;
 wire \u_delay_line.u_bulk_20.dl_4 ;
 wire \u_delay_line.u_bulk_20.dl_5 ;
 wire \u_delay_line.u_bulk_20.dl_6 ;
 wire \u_delay_line.u_bulk_20.dl_7 ;
 wire \u_delay_line.u_bulk_20.dl_8 ;
 wire \u_delay_line.u_bulk_20.dl_9 ;
 wire \u_delay_line.u_bulk_21.dl_0 ;
 wire \u_delay_line.u_bulk_21.dl_1 ;
 wire \u_delay_line.u_bulk_21.dl_10 ;
 wire \u_delay_line.u_bulk_21.dl_11 ;
 wire \u_delay_line.u_bulk_21.dl_12 ;
 wire \u_delay_line.u_bulk_21.dl_13 ;
 wire \u_delay_line.u_bulk_21.dl_14 ;
 wire \u_delay_line.u_bulk_21.dl_2 ;
 wire \u_delay_line.u_bulk_21.dl_3 ;
 wire \u_delay_line.u_bulk_21.dl_4 ;
 wire \u_delay_line.u_bulk_21.dl_5 ;
 wire \u_delay_line.u_bulk_21.dl_6 ;
 wire \u_delay_line.u_bulk_21.dl_7 ;
 wire \u_delay_line.u_bulk_21.dl_8 ;
 wire \u_delay_line.u_bulk_21.dl_9 ;
 wire \u_delay_line.u_bulk_3.dl_0 ;
 wire \u_delay_line.u_bulk_3.dl_1 ;
 wire \u_delay_line.u_bulk_3.dl_10 ;
 wire \u_delay_line.u_bulk_3.dl_11 ;
 wire \u_delay_line.u_bulk_3.dl_12 ;
 wire \u_delay_line.u_bulk_3.dl_13 ;
 wire \u_delay_line.u_bulk_3.dl_14 ;
 wire \u_delay_line.u_bulk_3.dl_2 ;
 wire \u_delay_line.u_bulk_3.dl_3 ;
 wire \u_delay_line.u_bulk_3.dl_4 ;
 wire \u_delay_line.u_bulk_3.dl_5 ;
 wire \u_delay_line.u_bulk_3.dl_6 ;
 wire \u_delay_line.u_bulk_3.dl_7 ;
 wire \u_delay_line.u_bulk_3.dl_8 ;
 wire \u_delay_line.u_bulk_3.dl_9 ;
 wire \u_delay_line.u_bulk_4.dl_0 ;
 wire \u_delay_line.u_bulk_4.dl_1 ;
 wire \u_delay_line.u_bulk_4.dl_10 ;
 wire \u_delay_line.u_bulk_4.dl_11 ;
 wire \u_delay_line.u_bulk_4.dl_12 ;
 wire \u_delay_line.u_bulk_4.dl_13 ;
 wire \u_delay_line.u_bulk_4.dl_14 ;
 wire \u_delay_line.u_bulk_4.dl_2 ;
 wire \u_delay_line.u_bulk_4.dl_3 ;
 wire \u_delay_line.u_bulk_4.dl_4 ;
 wire \u_delay_line.u_bulk_4.dl_5 ;
 wire \u_delay_line.u_bulk_4.dl_6 ;
 wire \u_delay_line.u_bulk_4.dl_7 ;
 wire \u_delay_line.u_bulk_4.dl_8 ;
 wire \u_delay_line.u_bulk_4.dl_9 ;
 wire \u_delay_line.u_bulk_5.dl_0 ;
 wire \u_delay_line.u_bulk_5.dl_1 ;
 wire \u_delay_line.u_bulk_5.dl_10 ;
 wire \u_delay_line.u_bulk_5.dl_11 ;
 wire \u_delay_line.u_bulk_5.dl_12 ;
 wire \u_delay_line.u_bulk_5.dl_13 ;
 wire \u_delay_line.u_bulk_5.dl_14 ;
 wire \u_delay_line.u_bulk_5.dl_2 ;
 wire \u_delay_line.u_bulk_5.dl_3 ;
 wire \u_delay_line.u_bulk_5.dl_4 ;
 wire \u_delay_line.u_bulk_5.dl_5 ;
 wire \u_delay_line.u_bulk_5.dl_6 ;
 wire \u_delay_line.u_bulk_5.dl_7 ;
 wire \u_delay_line.u_bulk_5.dl_8 ;
 wire \u_delay_line.u_bulk_5.dl_9 ;
 wire \u_delay_line.u_bulk_6.dl_0 ;
 wire \u_delay_line.u_bulk_6.dl_1 ;
 wire \u_delay_line.u_bulk_6.dl_10 ;
 wire \u_delay_line.u_bulk_6.dl_11 ;
 wire \u_delay_line.u_bulk_6.dl_12 ;
 wire \u_delay_line.u_bulk_6.dl_13 ;
 wire \u_delay_line.u_bulk_6.dl_14 ;
 wire \u_delay_line.u_bulk_6.dl_2 ;
 wire \u_delay_line.u_bulk_6.dl_3 ;
 wire \u_delay_line.u_bulk_6.dl_4 ;
 wire \u_delay_line.u_bulk_6.dl_5 ;
 wire \u_delay_line.u_bulk_6.dl_6 ;
 wire \u_delay_line.u_bulk_6.dl_7 ;
 wire \u_delay_line.u_bulk_6.dl_8 ;
 wire \u_delay_line.u_bulk_6.dl_9 ;
 wire \u_delay_line.u_bulk_7.dl_0 ;
 wire \u_delay_line.u_bulk_7.dl_1 ;
 wire \u_delay_line.u_bulk_7.dl_10 ;
 wire \u_delay_line.u_bulk_7.dl_11 ;
 wire \u_delay_line.u_bulk_7.dl_12 ;
 wire \u_delay_line.u_bulk_7.dl_13 ;
 wire \u_delay_line.u_bulk_7.dl_14 ;
 wire \u_delay_line.u_bulk_7.dl_2 ;
 wire \u_delay_line.u_bulk_7.dl_3 ;
 wire \u_delay_line.u_bulk_7.dl_4 ;
 wire \u_delay_line.u_bulk_7.dl_5 ;
 wire \u_delay_line.u_bulk_7.dl_6 ;
 wire \u_delay_line.u_bulk_7.dl_7 ;
 wire \u_delay_line.u_bulk_7.dl_8 ;
 wire \u_delay_line.u_bulk_7.dl_9 ;
 wire \u_delay_line.u_bulk_8.dl_0 ;
 wire \u_delay_line.u_bulk_8.dl_1 ;
 wire \u_delay_line.u_bulk_8.dl_10 ;
 wire \u_delay_line.u_bulk_8.dl_11 ;
 wire \u_delay_line.u_bulk_8.dl_12 ;
 wire \u_delay_line.u_bulk_8.dl_13 ;
 wire \u_delay_line.u_bulk_8.dl_14 ;
 wire \u_delay_line.u_bulk_8.dl_2 ;
 wire \u_delay_line.u_bulk_8.dl_3 ;
 wire \u_delay_line.u_bulk_8.dl_4 ;
 wire \u_delay_line.u_bulk_8.dl_5 ;
 wire \u_delay_line.u_bulk_8.dl_6 ;
 wire \u_delay_line.u_bulk_8.dl_7 ;
 wire \u_delay_line.u_bulk_8.dl_8 ;
 wire \u_delay_line.u_bulk_8.dl_9 ;
 wire \u_delay_line.u_bulk_9.dl_0 ;
 wire \u_delay_line.u_bulk_9.dl_1 ;
 wire \u_delay_line.u_bulk_9.dl_10 ;
 wire \u_delay_line.u_bulk_9.dl_11 ;
 wire \u_delay_line.u_bulk_9.dl_12 ;
 wire \u_delay_line.u_bulk_9.dl_13 ;
 wire \u_delay_line.u_bulk_9.dl_14 ;
 wire \u_delay_line.u_bulk_9.dl_2 ;
 wire \u_delay_line.u_bulk_9.dl_3 ;
 wire \u_delay_line.u_bulk_9.dl_4 ;
 wire \u_delay_line.u_bulk_9.dl_5 ;
 wire \u_delay_line.u_bulk_9.dl_6 ;
 wire \u_delay_line.u_bulk_9.dl_7 ;
 wire \u_delay_line.u_bulk_9.dl_8 ;
 wire \u_delay_line.u_bulk_9.dl_9 ;
 wire \u_delay_line.u_dl_0.dl_0 ;
 wire \u_delay_line.u_dl_0.dl_1 ;
 wire \u_delay_line.u_dl_0.dl_10 ;
 wire \u_delay_line.u_dl_0.dl_2 ;
 wire \u_delay_line.u_dl_0.dl_3 ;
 wire \u_delay_line.u_dl_0.dl_4 ;
 wire \u_delay_line.u_dl_0.dl_5 ;
 wire \u_delay_line.u_dl_0.dl_6 ;
 wire \u_delay_line.u_dl_0.dl_7 ;
 wire \u_delay_line.u_dl_0.dl_8 ;
 wire \u_delay_line.u_dl_0.dl_9 ;
 wire \u_delay_line.u_dl_1.dl_0 ;
 wire \u_delay_line.u_dl_1.dl_1 ;
 wire \u_delay_line.u_dl_1.dl_10 ;
 wire \u_delay_line.u_dl_1.dl_2 ;
 wire \u_delay_line.u_dl_1.dl_3 ;
 wire \u_delay_line.u_dl_1.dl_4 ;
 wire \u_delay_line.u_dl_1.dl_5 ;
 wire \u_delay_line.u_dl_1.dl_6 ;
 wire \u_delay_line.u_dl_1.dl_7 ;
 wire \u_delay_line.u_dl_1.dl_8 ;
 wire \u_delay_line.u_dl_1.dl_9 ;
 wire \u_delay_line.u_dl_10.dl_0 ;
 wire \u_delay_line.u_dl_10.dl_1 ;
 wire \u_delay_line.u_dl_10.dl_10 ;
 wire \u_delay_line.u_dl_10.dl_2 ;
 wire \u_delay_line.u_dl_10.dl_3 ;
 wire \u_delay_line.u_dl_10.dl_4 ;
 wire \u_delay_line.u_dl_10.dl_5 ;
 wire \u_delay_line.u_dl_10.dl_6 ;
 wire \u_delay_line.u_dl_10.dl_7 ;
 wire \u_delay_line.u_dl_10.dl_8 ;
 wire \u_delay_line.u_dl_10.dl_9 ;
 wire \u_delay_line.u_dl_11.dl_0 ;
 wire \u_delay_line.u_dl_11.dl_1 ;
 wire \u_delay_line.u_dl_11.dl_10 ;
 wire \u_delay_line.u_dl_11.dl_2 ;
 wire \u_delay_line.u_dl_11.dl_3 ;
 wire \u_delay_line.u_dl_11.dl_4 ;
 wire \u_delay_line.u_dl_11.dl_5 ;
 wire \u_delay_line.u_dl_11.dl_6 ;
 wire \u_delay_line.u_dl_11.dl_7 ;
 wire \u_delay_line.u_dl_11.dl_8 ;
 wire \u_delay_line.u_dl_11.dl_9 ;
 wire \u_delay_line.u_dl_12.dl_0 ;
 wire \u_delay_line.u_dl_12.dl_1 ;
 wire \u_delay_line.u_dl_12.dl_10 ;
 wire \u_delay_line.u_dl_12.dl_2 ;
 wire \u_delay_line.u_dl_12.dl_3 ;
 wire \u_delay_line.u_dl_12.dl_4 ;
 wire \u_delay_line.u_dl_12.dl_5 ;
 wire \u_delay_line.u_dl_12.dl_6 ;
 wire \u_delay_line.u_dl_12.dl_7 ;
 wire \u_delay_line.u_dl_12.dl_8 ;
 wire \u_delay_line.u_dl_12.dl_9 ;
 wire \u_delay_line.u_dl_13.dl_0 ;
 wire \u_delay_line.u_dl_13.dl_1 ;
 wire \u_delay_line.u_dl_13.dl_10 ;
 wire \u_delay_line.u_dl_13.dl_2 ;
 wire \u_delay_line.u_dl_13.dl_3 ;
 wire \u_delay_line.u_dl_13.dl_4 ;
 wire \u_delay_line.u_dl_13.dl_5 ;
 wire \u_delay_line.u_dl_13.dl_6 ;
 wire \u_delay_line.u_dl_13.dl_7 ;
 wire \u_delay_line.u_dl_13.dl_8 ;
 wire \u_delay_line.u_dl_13.dl_9 ;
 wire \u_delay_line.u_dl_14.dl_0 ;
 wire \u_delay_line.u_dl_14.dl_1 ;
 wire \u_delay_line.u_dl_14.dl_10 ;
 wire \u_delay_line.u_dl_14.dl_2 ;
 wire \u_delay_line.u_dl_14.dl_3 ;
 wire \u_delay_line.u_dl_14.dl_4 ;
 wire \u_delay_line.u_dl_14.dl_5 ;
 wire \u_delay_line.u_dl_14.dl_6 ;
 wire \u_delay_line.u_dl_14.dl_7 ;
 wire \u_delay_line.u_dl_14.dl_8 ;
 wire \u_delay_line.u_dl_14.dl_9 ;
 wire \u_delay_line.u_dl_15.dl_0 ;
 wire \u_delay_line.u_dl_15.dl_1 ;
 wire \u_delay_line.u_dl_15.dl_10 ;
 wire \u_delay_line.u_dl_15.dl_2 ;
 wire \u_delay_line.u_dl_15.dl_3 ;
 wire \u_delay_line.u_dl_15.dl_4 ;
 wire \u_delay_line.u_dl_15.dl_5 ;
 wire \u_delay_line.u_dl_15.dl_6 ;
 wire \u_delay_line.u_dl_15.dl_7 ;
 wire \u_delay_line.u_dl_15.dl_8 ;
 wire \u_delay_line.u_dl_15.dl_9 ;
 wire \u_delay_line.u_dl_16.dl_0 ;
 wire \u_delay_line.u_dl_16.dl_1 ;
 wire \u_delay_line.u_dl_16.dl_10 ;
 wire \u_delay_line.u_dl_16.dl_2 ;
 wire \u_delay_line.u_dl_16.dl_3 ;
 wire \u_delay_line.u_dl_16.dl_4 ;
 wire \u_delay_line.u_dl_16.dl_5 ;
 wire \u_delay_line.u_dl_16.dl_6 ;
 wire \u_delay_line.u_dl_16.dl_7 ;
 wire \u_delay_line.u_dl_16.dl_8 ;
 wire \u_delay_line.u_dl_16.dl_9 ;
 wire \u_delay_line.u_dl_17.dl_0 ;
 wire \u_delay_line.u_dl_17.dl_1 ;
 wire \u_delay_line.u_dl_17.dl_10 ;
 wire \u_delay_line.u_dl_17.dl_2 ;
 wire \u_delay_line.u_dl_17.dl_3 ;
 wire \u_delay_line.u_dl_17.dl_4 ;
 wire \u_delay_line.u_dl_17.dl_5 ;
 wire \u_delay_line.u_dl_17.dl_6 ;
 wire \u_delay_line.u_dl_17.dl_7 ;
 wire \u_delay_line.u_dl_17.dl_8 ;
 wire \u_delay_line.u_dl_17.dl_9 ;
 wire \u_delay_line.u_dl_18.dl_0 ;
 wire \u_delay_line.u_dl_18.dl_1 ;
 wire \u_delay_line.u_dl_18.dl_10 ;
 wire \u_delay_line.u_dl_18.dl_2 ;
 wire \u_delay_line.u_dl_18.dl_3 ;
 wire \u_delay_line.u_dl_18.dl_4 ;
 wire \u_delay_line.u_dl_18.dl_5 ;
 wire \u_delay_line.u_dl_18.dl_6 ;
 wire \u_delay_line.u_dl_18.dl_7 ;
 wire \u_delay_line.u_dl_18.dl_8 ;
 wire \u_delay_line.u_dl_18.dl_9 ;
 wire \u_delay_line.u_dl_19.dl_0 ;
 wire \u_delay_line.u_dl_19.dl_1 ;
 wire \u_delay_line.u_dl_19.dl_10 ;
 wire \u_delay_line.u_dl_19.dl_2 ;
 wire \u_delay_line.u_dl_19.dl_3 ;
 wire \u_delay_line.u_dl_19.dl_4 ;
 wire \u_delay_line.u_dl_19.dl_5 ;
 wire \u_delay_line.u_dl_19.dl_6 ;
 wire \u_delay_line.u_dl_19.dl_7 ;
 wire \u_delay_line.u_dl_19.dl_8 ;
 wire \u_delay_line.u_dl_19.dl_9 ;
 wire \u_delay_line.u_dl_2.dl_0 ;
 wire \u_delay_line.u_dl_2.dl_1 ;
 wire \u_delay_line.u_dl_2.dl_10 ;
 wire \u_delay_line.u_dl_2.dl_2 ;
 wire \u_delay_line.u_dl_2.dl_3 ;
 wire \u_delay_line.u_dl_2.dl_4 ;
 wire \u_delay_line.u_dl_2.dl_5 ;
 wire \u_delay_line.u_dl_2.dl_6 ;
 wire \u_delay_line.u_dl_2.dl_7 ;
 wire \u_delay_line.u_dl_2.dl_8 ;
 wire \u_delay_line.u_dl_2.dl_9 ;
 wire \u_delay_line.u_dl_20.dl_0 ;
 wire \u_delay_line.u_dl_20.dl_1 ;
 wire \u_delay_line.u_dl_20.dl_10 ;
 wire \u_delay_line.u_dl_20.dl_2 ;
 wire \u_delay_line.u_dl_20.dl_3 ;
 wire \u_delay_line.u_dl_20.dl_4 ;
 wire \u_delay_line.u_dl_20.dl_5 ;
 wire \u_delay_line.u_dl_20.dl_6 ;
 wire \u_delay_line.u_dl_20.dl_7 ;
 wire \u_delay_line.u_dl_20.dl_8 ;
 wire \u_delay_line.u_dl_20.dl_9 ;
 wire \u_delay_line.u_dl_21.dl_0 ;
 wire \u_delay_line.u_dl_21.dl_1 ;
 wire \u_delay_line.u_dl_21.dl_10 ;
 wire \u_delay_line.u_dl_21.dl_2 ;
 wire \u_delay_line.u_dl_21.dl_3 ;
 wire \u_delay_line.u_dl_21.dl_4 ;
 wire \u_delay_line.u_dl_21.dl_5 ;
 wire \u_delay_line.u_dl_21.dl_6 ;
 wire \u_delay_line.u_dl_21.dl_7 ;
 wire \u_delay_line.u_dl_21.dl_8 ;
 wire \u_delay_line.u_dl_21.dl_9 ;
 wire \u_delay_line.u_dl_22.dl_0 ;
 wire \u_delay_line.u_dl_22.dl_1 ;
 wire \u_delay_line.u_dl_22.dl_10 ;
 wire \u_delay_line.u_dl_22.dl_2 ;
 wire \u_delay_line.u_dl_22.dl_3 ;
 wire \u_delay_line.u_dl_22.dl_4 ;
 wire \u_delay_line.u_dl_22.dl_5 ;
 wire \u_delay_line.u_dl_22.dl_6 ;
 wire \u_delay_line.u_dl_22.dl_7 ;
 wire \u_delay_line.u_dl_22.dl_8 ;
 wire \u_delay_line.u_dl_22.dl_9 ;
 wire \u_delay_line.u_dl_23.dl_0 ;
 wire \u_delay_line.u_dl_23.dl_1 ;
 wire \u_delay_line.u_dl_23.dl_10 ;
 wire \u_delay_line.u_dl_23.dl_2 ;
 wire \u_delay_line.u_dl_23.dl_3 ;
 wire \u_delay_line.u_dl_23.dl_4 ;
 wire \u_delay_line.u_dl_23.dl_5 ;
 wire \u_delay_line.u_dl_23.dl_6 ;
 wire \u_delay_line.u_dl_23.dl_7 ;
 wire \u_delay_line.u_dl_23.dl_8 ;
 wire \u_delay_line.u_dl_23.dl_9 ;
 wire \u_delay_line.u_dl_24.dl_0 ;
 wire \u_delay_line.u_dl_24.dl_1 ;
 wire \u_delay_line.u_dl_24.dl_10 ;
 wire \u_delay_line.u_dl_24.dl_2 ;
 wire \u_delay_line.u_dl_24.dl_3 ;
 wire \u_delay_line.u_dl_24.dl_4 ;
 wire \u_delay_line.u_dl_24.dl_5 ;
 wire \u_delay_line.u_dl_24.dl_6 ;
 wire \u_delay_line.u_dl_24.dl_7 ;
 wire \u_delay_line.u_dl_24.dl_8 ;
 wire \u_delay_line.u_dl_24.dl_9 ;
 wire \u_delay_line.u_dl_25.dl_0 ;
 wire \u_delay_line.u_dl_25.dl_1 ;
 wire \u_delay_line.u_dl_25.dl_10 ;
 wire \u_delay_line.u_dl_25.dl_2 ;
 wire \u_delay_line.u_dl_25.dl_3 ;
 wire \u_delay_line.u_dl_25.dl_4 ;
 wire \u_delay_line.u_dl_25.dl_5 ;
 wire \u_delay_line.u_dl_25.dl_6 ;
 wire \u_delay_line.u_dl_25.dl_7 ;
 wire \u_delay_line.u_dl_25.dl_8 ;
 wire \u_delay_line.u_dl_25.dl_9 ;
 wire \u_delay_line.u_dl_26.dl_0 ;
 wire \u_delay_line.u_dl_26.dl_1 ;
 wire \u_delay_line.u_dl_26.dl_10 ;
 wire \u_delay_line.u_dl_26.dl_2 ;
 wire \u_delay_line.u_dl_26.dl_3 ;
 wire \u_delay_line.u_dl_26.dl_4 ;
 wire \u_delay_line.u_dl_26.dl_5 ;
 wire \u_delay_line.u_dl_26.dl_6 ;
 wire \u_delay_line.u_dl_26.dl_7 ;
 wire \u_delay_line.u_dl_26.dl_8 ;
 wire \u_delay_line.u_dl_26.dl_9 ;
 wire \u_delay_line.u_dl_27.dl_0 ;
 wire \u_delay_line.u_dl_27.dl_1 ;
 wire \u_delay_line.u_dl_27.dl_10 ;
 wire \u_delay_line.u_dl_27.dl_2 ;
 wire \u_delay_line.u_dl_27.dl_3 ;
 wire \u_delay_line.u_dl_27.dl_4 ;
 wire \u_delay_line.u_dl_27.dl_5 ;
 wire \u_delay_line.u_dl_27.dl_6 ;
 wire \u_delay_line.u_dl_27.dl_7 ;
 wire \u_delay_line.u_dl_27.dl_8 ;
 wire \u_delay_line.u_dl_27.dl_9 ;
 wire \u_delay_line.u_dl_28.dl_0 ;
 wire \u_delay_line.u_dl_28.dl_1 ;
 wire \u_delay_line.u_dl_28.dl_10 ;
 wire \u_delay_line.u_dl_28.dl_2 ;
 wire \u_delay_line.u_dl_28.dl_3 ;
 wire \u_delay_line.u_dl_28.dl_4 ;
 wire \u_delay_line.u_dl_28.dl_5 ;
 wire \u_delay_line.u_dl_28.dl_6 ;
 wire \u_delay_line.u_dl_28.dl_7 ;
 wire \u_delay_line.u_dl_28.dl_8 ;
 wire \u_delay_line.u_dl_28.dl_9 ;
 wire \u_delay_line.u_dl_29.dl_0 ;
 wire \u_delay_line.u_dl_29.dl_1 ;
 wire \u_delay_line.u_dl_29.dl_10 ;
 wire \u_delay_line.u_dl_29.dl_2 ;
 wire \u_delay_line.u_dl_29.dl_3 ;
 wire \u_delay_line.u_dl_29.dl_4 ;
 wire \u_delay_line.u_dl_29.dl_5 ;
 wire \u_delay_line.u_dl_29.dl_6 ;
 wire \u_delay_line.u_dl_29.dl_7 ;
 wire \u_delay_line.u_dl_29.dl_8 ;
 wire \u_delay_line.u_dl_29.dl_9 ;
 wire \u_delay_line.u_dl_3.dl_0 ;
 wire \u_delay_line.u_dl_3.dl_1 ;
 wire \u_delay_line.u_dl_3.dl_10 ;
 wire \u_delay_line.u_dl_3.dl_2 ;
 wire \u_delay_line.u_dl_3.dl_3 ;
 wire \u_delay_line.u_dl_3.dl_4 ;
 wire \u_delay_line.u_dl_3.dl_5 ;
 wire \u_delay_line.u_dl_3.dl_6 ;
 wire \u_delay_line.u_dl_3.dl_7 ;
 wire \u_delay_line.u_dl_3.dl_8 ;
 wire \u_delay_line.u_dl_3.dl_9 ;
 wire \u_delay_line.u_dl_30.dl_0 ;
 wire \u_delay_line.u_dl_30.dl_1 ;
 wire \u_delay_line.u_dl_30.dl_10 ;
 wire \u_delay_line.u_dl_30.dl_2 ;
 wire \u_delay_line.u_dl_30.dl_3 ;
 wire \u_delay_line.u_dl_30.dl_4 ;
 wire \u_delay_line.u_dl_30.dl_5 ;
 wire \u_delay_line.u_dl_30.dl_6 ;
 wire \u_delay_line.u_dl_30.dl_7 ;
 wire \u_delay_line.u_dl_30.dl_8 ;
 wire \u_delay_line.u_dl_30.dl_9 ;
 wire \u_delay_line.u_dl_31.dl_0 ;
 wire \u_delay_line.u_dl_31.dl_1 ;
 wire \u_delay_line.u_dl_31.dl_10 ;
 wire \u_delay_line.u_dl_31.dl_2 ;
 wire \u_delay_line.u_dl_31.dl_3 ;
 wire \u_delay_line.u_dl_31.dl_4 ;
 wire \u_delay_line.u_dl_31.dl_5 ;
 wire \u_delay_line.u_dl_31.dl_6 ;
 wire \u_delay_line.u_dl_31.dl_7 ;
 wire \u_delay_line.u_dl_31.dl_8 ;
 wire \u_delay_line.u_dl_31.dl_9 ;
 wire \u_delay_line.u_dl_4.dl_0 ;
 wire \u_delay_line.u_dl_4.dl_1 ;
 wire \u_delay_line.u_dl_4.dl_10 ;
 wire \u_delay_line.u_dl_4.dl_2 ;
 wire \u_delay_line.u_dl_4.dl_3 ;
 wire \u_delay_line.u_dl_4.dl_4 ;
 wire \u_delay_line.u_dl_4.dl_5 ;
 wire \u_delay_line.u_dl_4.dl_6 ;
 wire \u_delay_line.u_dl_4.dl_7 ;
 wire \u_delay_line.u_dl_4.dl_8 ;
 wire \u_delay_line.u_dl_4.dl_9 ;
 wire \u_delay_line.u_dl_5.dl_0 ;
 wire \u_delay_line.u_dl_5.dl_1 ;
 wire \u_delay_line.u_dl_5.dl_10 ;
 wire \u_delay_line.u_dl_5.dl_2 ;
 wire \u_delay_line.u_dl_5.dl_3 ;
 wire \u_delay_line.u_dl_5.dl_4 ;
 wire \u_delay_line.u_dl_5.dl_5 ;
 wire \u_delay_line.u_dl_5.dl_6 ;
 wire \u_delay_line.u_dl_5.dl_7 ;
 wire \u_delay_line.u_dl_5.dl_8 ;
 wire \u_delay_line.u_dl_5.dl_9 ;
 wire \u_delay_line.u_dl_6.dl_0 ;
 wire \u_delay_line.u_dl_6.dl_1 ;
 wire \u_delay_line.u_dl_6.dl_10 ;
 wire \u_delay_line.u_dl_6.dl_2 ;
 wire \u_delay_line.u_dl_6.dl_3 ;
 wire \u_delay_line.u_dl_6.dl_4 ;
 wire \u_delay_line.u_dl_6.dl_5 ;
 wire \u_delay_line.u_dl_6.dl_6 ;
 wire \u_delay_line.u_dl_6.dl_7 ;
 wire \u_delay_line.u_dl_6.dl_8 ;
 wire \u_delay_line.u_dl_6.dl_9 ;
 wire \u_delay_line.u_dl_7.dl_0 ;
 wire \u_delay_line.u_dl_7.dl_1 ;
 wire \u_delay_line.u_dl_7.dl_10 ;
 wire \u_delay_line.u_dl_7.dl_2 ;
 wire \u_delay_line.u_dl_7.dl_3 ;
 wire \u_delay_line.u_dl_7.dl_4 ;
 wire \u_delay_line.u_dl_7.dl_5 ;
 wire \u_delay_line.u_dl_7.dl_6 ;
 wire \u_delay_line.u_dl_7.dl_7 ;
 wire \u_delay_line.u_dl_7.dl_8 ;
 wire \u_delay_line.u_dl_7.dl_9 ;
 wire \u_delay_line.u_dl_8.dl_0 ;
 wire \u_delay_line.u_dl_8.dl_1 ;
 wire \u_delay_line.u_dl_8.dl_10 ;
 wire \u_delay_line.u_dl_8.dl_2 ;
 wire \u_delay_line.u_dl_8.dl_3 ;
 wire \u_delay_line.u_dl_8.dl_4 ;
 wire \u_delay_line.u_dl_8.dl_5 ;
 wire \u_delay_line.u_dl_8.dl_6 ;
 wire \u_delay_line.u_dl_8.dl_7 ;
 wire \u_delay_line.u_dl_8.dl_8 ;
 wire \u_delay_line.u_dl_8.dl_9 ;
 wire \u_delay_line.u_dl_9.dl_0 ;
 wire \u_delay_line.u_dl_9.dl_1 ;
 wire \u_delay_line.u_dl_9.dl_10 ;
 wire \u_delay_line.u_dl_9.dl_2 ;
 wire \u_delay_line.u_dl_9.dl_3 ;
 wire \u_delay_line.u_dl_9.dl_4 ;
 wire \u_delay_line.u_dl_9.dl_5 ;
 wire \u_delay_line.u_dl_9.dl_6 ;
 wire \u_delay_line.u_dl_9.dl_7 ;
 wire \u_delay_line.u_dl_9.dl_8 ;
 wire \u_delay_line.u_dl_9.dl_9 ;
 wire \u_delay_line.valid_d ;
 wire \u_delay_line.valid_q ;
 wire \u_driver.data_dl[32] ;
 wire \u_driver.data_dl[33] ;
 wire \u_driver.data_dl[34] ;
 wire \u_driver.data_dl[35] ;
 wire \u_driver.data_dl[36] ;
 wire \u_driver.data_dl[37] ;
 wire \u_driver.data_dl[38] ;
 wire \u_driver.data_dl[39] ;
 wire \u_driver.data_edge[13] ;
 wire \u_driver.data_edge[14] ;
 wire \u_driver.data_edge[15] ;
 wire \u_driver.data_edge[16] ;
 wire \u_driver.data_edge[17] ;
 wire \u_driver.data_edge[18] ;
 wire \u_driver.data_edge[19] ;
 wire \u_driver.data_edge[20] ;
 wire \u_driver.data_edge[21] ;
 wire \u_driver.data_edge[22] ;
 wire \u_driver.data_edge[23] ;
 wire \u_driver.data_edge[24] ;
 wire \u_driver.data_edge[25] ;
 wire \u_driver.data_edge[26] ;
 wire \u_driver.data_edge[27] ;
 wire \u_driver.data_edge[28] ;
 wire \u_driver.data_edge[29] ;
 wire \u_driver.data_edge[30] ;
 wire \u_driver.data_edge[31] ;
 wire \u_driver.data_edge[32] ;
 wire \u_driver.data_edge[33] ;
 wire \u_driver.data_edge[34] ;
 wire \u_driver.data_edge[35] ;
 wire \u_driver.data_edge[36] ;
 wire \u_driver.data_edge[37] ;
 wire \u_driver.data_edge[38] ;
 wire \u_driver.data_edge[39] ;
 wire \u_driver.data_in[0] ;
 wire \u_driver.data_in[1] ;
 wire \u_driver.data_in[2] ;
 wire \u_driver.data_in[39] ;
 wire \u_driver.data_in[3] ;
 wire \u_driver.data_q[36] ;
 wire \u_driver.data_q[37] ;
 wire \u_driver.data_q[38] ;
 wire \u_driver.data_q[39] ;
 wire \u_driver.dl_en ;
 wire \u_driver.edge_cnt_q[0] ;
 wire \u_driver.edge_cnt_q[1] ;
 wire \u_driver.edge_cnt_q[2] ;
 wire \u_driver.edge_cnt_q[3] ;
 wire \u_driver.i_data[0] ;
 wire \u_driver.i_data[1] ;
 wire \u_driver.i_data[2] ;
 wire \u_driver.i_data[3] ;
 wire \u_driver.i_valid ;
 wire \u_driver.o_valid ;
 wire \u_driver.p1_capture ;
 wire \u_rx.p1_rx ;
 wire \u_rx.sm_uart_q[0] ;
 wire \u_rx.sm_uart_q[1] ;
 wire \u_rx.sm_uart_q[2] ;
 wire \u_rx.sm_uart_q[3] ;
 wire \u_rx.timer_q[0] ;
 wire \u_rx.timer_q[10] ;
 wire \u_rx.timer_q[11] ;
 wire \u_rx.timer_q[12] ;
 wire \u_rx.timer_q[1] ;
 wire \u_rx.timer_q[2] ;
 wire \u_rx.timer_q[3] ;
 wire \u_rx.timer_q[4] ;
 wire \u_rx.timer_q[5] ;
 wire \u_rx.timer_q[6] ;
 wire \u_rx.timer_q[7] ;
 wire \u_rx.timer_q[8] ;
 wire \u_rx.timer_q[9] ;
 wire \u_rx.valid_d ;
 wire \u_tx.o_tx ;
 wire \u_tx.sm_uart_q[0] ;
 wire \u_tx.sm_uart_q[1] ;
 wire \u_tx.sm_uart_q[2] ;
 wire \u_tx.sm_uart_q[3] ;
 wire \u_tx.sm_uart_q[4] ;
 wire \u_tx.timer_q[0] ;
 wire \u_tx.timer_q[10] ;
 wire \u_tx.timer_q[11] ;
 wire \u_tx.timer_q[12] ;
 wire \u_tx.timer_q[1] ;
 wire \u_tx.timer_q[2] ;
 wire \u_tx.timer_q[3] ;
 wire \u_tx.timer_q[4] ;
 wire \u_tx.timer_q[5] ;
 wire \u_tx.timer_q[6] ;
 wire \u_tx.timer_q[7] ;
 wire \u_tx.timer_q[8] ;
 wire \u_tx.timer_q[9] ;

 sky130_fd_sc_hd__decap_8 FILLER_0_0_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_121 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_0_134 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_144 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_0_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_156 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_176 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_184 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_209 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_221 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_256 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_260 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_264 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_277 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_0_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_289 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_298 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_0_32 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_337 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_349 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_38 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_0_64 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_70 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_0_91 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_99 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_10_119 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_123 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_134 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_10_18 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_10_192 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_205 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_10_237 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_241 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_10_268 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_10_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_295 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_10_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_329 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_33 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_350 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_60 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_10_67 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_71 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_10_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_91 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_104 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_11_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_119 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_146 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_11_158 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_11_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_11_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_11_17 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_175 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_11_184 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_190 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_211 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_11_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_231 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_243 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_11_25 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_264 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_11_276 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_11_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_285 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_11_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_321 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_11_329 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_335 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_11_345 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_40 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_11_52 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_11_64 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_11_92 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_11_98 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_115 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_124 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_12_136 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_12_157 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_12_16 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_12_189 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_12_205 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_211 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_12_219 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_12_233 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_24 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_12_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_257 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_270 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_12_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_12_305 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_312 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_350 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_12_78 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_12_91 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_99 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_13_104 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_13_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_117 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_13_12 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_13_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_13_150 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_13_156 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_178 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_13_190 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_13_221 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_13_252 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_13_270 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_13_275 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_13_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_301 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_313 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_13_325 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_33 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_13_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_337 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_13_349 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_13_45 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_13_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_13_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_13_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_13_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_103 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_14_112 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_14_132 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_14_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_147 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_14_152 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_158 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_14_165 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_176 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_14_185 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_14_193 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_205 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_14_224 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_239 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_14_247 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_14_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_259 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_266 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_278 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_290 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_14_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_14_302 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_14_32 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_14_349 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_40 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_47 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_71 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_14_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_91 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_101 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_15_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_117 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_15_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_157 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_15_165 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_15_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_179 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_15_18 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_188 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_15_220 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_237 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_15_254 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_270 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_15_274 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_15_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_301 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_15_31 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_15_316 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_320 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_15_329 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_335 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_349 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_45 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_15_72 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_76 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_15_94 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_121 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_16_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_16_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_16_154 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_16_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_174 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_16_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_16_190 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_16_218 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_238 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_16_248 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_16_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_272 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_293 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_16_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_16_305 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_315 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_16_32 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_16_320 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_349 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_36 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_46 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_16_91 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_99 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_17_107 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_17_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_17_126 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_17_134 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_14 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_17_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_17_179 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_17_203 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_214 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_17_254 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_262 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_17_269 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_17_277 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_17_293 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_299 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_17_324 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_17_337 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_17_346 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_350 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_17_36 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_17_45 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_17_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_17_70 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_17_78 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_95 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_18_112 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_18_134 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_18_147 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_18_163 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_18_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_18_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_18_221 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_18_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_266 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_18_290 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_18_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_18_301 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_18_321 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_18_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_50 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_56 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_18_68 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_76 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_92 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_19_108 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_19_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_19_146 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_19_16 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_19_164 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_176 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_19_216 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_19_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_19_234 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_243 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_19_255 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_267 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_293 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_19_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_19_308 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_19_316 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_19_322 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_326 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_335 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_19_337 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_341 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_19_346 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_350 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_19_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_19_75 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_87 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_99 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_1_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_1_119 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_1_148 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_1_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_1_175 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_179 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_1_222 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_237 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_249 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_1_261 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_1_273 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_1_306 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_1_314 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_32 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_1_345 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_1_36 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_44 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_20_114 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_14 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_20_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_20_155 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_20_165 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_179 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_20_191 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_205 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_20_212 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_20_224 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_228 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_20_249 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_20_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_20_283 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_20_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_20_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_20_326 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_350 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_20_50 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_20_58 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_67 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_20_79 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_20_91 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_10 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_21_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_21_118 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_126 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_21_135 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_21_146 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_150 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_155 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_21_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_17 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_196 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_208 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_214 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_21_220 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_21_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_21_238 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_24 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_21_246 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_261 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_21_273 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_21_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_289 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_297 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_302 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_31 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_21_314 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_21_327 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_335 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_21_337 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_36 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_21_48 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_21_79 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_103 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_22_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_161 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_173 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_22_185 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_189 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_22_229 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_22_258 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_22_284 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_22_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_22_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_306 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_22_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_349 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_37 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_64 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_22_76 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_22_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_91 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_23_108 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_23_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_23_151 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_23_164 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_23_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_23_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_23_186 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_206 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_23_218 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_23_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_229 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_236 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_23_24 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_23_248 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_23_273 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_23_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_23_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_23_298 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_23_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_302 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_23_310 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_23_332 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_23_345 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_23_46 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_23_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_23_63 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_67 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_102 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_24_114 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_24_12 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_24_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_24_184 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_24_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_24_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_24_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_24_239 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_24_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_24_262 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_270 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_24_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_24_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_24_318 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_24_32 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_24_324 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_24_349 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_24_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_49 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_59 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_24_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_24_80 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_24_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_24_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_98 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_107 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_116 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_25_128 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_25_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_25_151 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_159 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_25_163 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_178 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_25_190 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_196 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_206 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_25_218 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_25_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_25_240 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_278 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_25_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_25_322 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_25_329 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_335 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_25_345 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_25_62 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_25_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_25_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_26_100 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_26_12 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_127 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_26_175 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_26_190 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_26_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_26_265 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_26_296 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_26_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_304 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_32 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_321 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_350 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_44 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_56 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_26_68 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_27_103 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_27_12 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_27_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_27_131 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_27_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_27_155 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_27_161 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_27_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_27_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_200 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_212 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_27_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_231 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_27_25 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_27_255 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_27_267 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_27_278 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_27_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_27_30 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_323 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_335 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_27_337 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_343 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_350 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_27_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_61 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_118 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_28_12 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_28_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_28_174 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_209 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_28_241 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_28_249 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_277 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_289 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_28_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_28_301 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_28_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_28_317 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_33 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_28_344 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_350 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_46 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_28_50 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_28_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_28_61 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_72 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_28_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_29_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_29_121 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_140 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_152 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_29_16 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_29_161 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_29_174 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_29_218 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_22 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_248 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_260 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_29_272 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_29_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_29_291 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_29_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_29_331 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_335 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_29_349 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_29_38 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_29_45 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_50 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_29_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_29_60 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_66 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_29_76 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_84 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_94 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_2_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_117 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_2_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_2_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_2_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_159 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_180 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_2_192 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_209 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_2_221 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_2_229 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_238 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_2_271 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_277 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_2_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_2_296 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_2_326 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_330 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_2_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_2_60 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_2_68 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_2_74 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_2_89 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_106 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_30_127 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_135 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_30_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_30_209 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_30_224 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_30_239 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_245 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_296 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_30_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_30_303 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_30_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_319 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_327 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_49 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_30_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_30_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_30_76 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_31_102 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_31_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_117 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_31_134 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_31_14 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_31_146 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_158 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_31_163 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_31_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_175 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_31_188 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_31_200 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_208 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_31_215 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_22 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_31_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_229 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_31_273 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_31_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_31_293 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_299 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_31_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_31_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_317 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_330 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_31_337 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_341 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_31_348 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_31_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_31_47 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_31_63 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_31_90 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_32_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_117 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_32_123 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_32_131 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_32_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_32_161 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_173 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_32_180 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_32_192 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_32_219 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_32_233 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_32_245 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_32_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_32_264 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_272 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_32_278 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_32_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_32_301 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_32_315 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_32_330 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_32_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_32_60 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_32_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_32_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_33_102 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_120 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_33_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_149 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_158 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_33_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_33_188 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_33_200 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_33_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_216 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_33_249 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_270 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_33_297 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_33_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_33_314 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_322 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_33 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_33_332 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_33_337 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_341 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_33_348 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_37 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_33_44 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_33_79 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_34_101 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_34_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_34_119 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_34_131 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_135 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_34_146 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_34_158 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_34_172 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_178 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_34_193 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_217 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_239 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_24 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_34_243 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_34_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_259 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_34_265 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_34_277 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_34_287 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_34_293 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_34_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_34_315 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_319 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_34_332 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_337 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_350 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_34_36 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_40 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_34_50 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_34_59 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_34_71 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_34_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_34_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_35_126 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_35_142 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_35_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_35_165 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_35_176 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_35_188 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_35_196 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_35_207 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_35_219 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_35_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_35_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_35_277 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_35_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_35_302 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_31 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_35_318 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_322 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_335 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_35_337 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_349 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_35_88 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_36_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_149 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_178 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_36_186 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_36_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_217 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_36_22 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_230 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_234 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_36_238 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_36_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_36_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_36_266 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_270 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_36_274 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_36_288 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_292 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_36_296 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_36_312 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_32 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_36_320 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_36_325 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_36_337 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_36_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_36_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_36_62 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_36_74 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_36_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_88 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_36_98 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_120 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_124 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_128 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_132 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_37_136 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_37_142 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_37_150 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_156 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_37_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_18 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_37_189 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_37_202 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_208 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_213 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_37_217 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_37_22 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_37_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_37_237 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_243 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_247 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_37_252 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_37_296 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_37_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_37_308 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_318 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_37_34 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_349 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_42 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_70 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_37_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_96 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_38_102 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_106 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_38_118 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_122 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_38_126 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_130 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_134 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_144 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_151 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_158 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_175 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_182 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_203 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_208 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_212 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_219 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_38_249 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_38_259 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_38_271 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_38_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_38_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_321 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_330 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_335 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_349 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_38 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_38_48 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_38_62 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_66 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_38_70 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_74 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_78 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_38_94 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_98 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_3_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_3_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_155 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_3_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_3_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_203 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_3_231 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_239 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_260 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_3_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_292 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_3_319 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_323 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_3_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_337 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_3_40 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_48 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_63 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_75 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_3_87 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_91 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_117 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_4_13 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_4_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_4_170 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_178 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_4_189 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_203 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_207 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_4_219 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_4_242 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_294 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_4_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_306 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_4_326 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_330 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_59 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_4_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_4_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_89 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_99 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_5_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_145 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_157 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_5_17 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_172 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_5_190 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_5_214 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_222 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_248 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_260 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_5_272 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_293 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_5_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_5_305 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_315 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_5_325 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_5_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_337 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_5_347 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_5_37 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_45 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_60 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_5_72 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_76 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_89 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_6_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_6_162 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_173 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_6_185 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_6_193 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_6_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_6_20 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_6_206 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_214 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_6_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_231 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_6_237 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_6_243 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_6_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_6_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_6_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_324 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_6_345 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_6_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_6_79 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_6_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_7_107 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_12 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_7_162 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_7_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_7_185 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_7_204 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_7_219 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_7_232 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_240 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_265 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_7_277 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_293 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_7_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_7_319 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_7_331 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_335 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_7_337 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_7_34 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_343 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_350 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_7_52 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_60 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_72 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_84 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_7_96 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_8_126 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_130 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_8_136 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_8_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_147 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_8_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_8_22 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_8_222 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_8_232 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_265 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_287 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_8_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_8_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_38 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_48 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_8_79 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_9_118 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_9_146 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_154 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_9_163 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_207 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_9_219 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_9_232 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_9_277 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_293 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_9_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_9_305 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_9_315 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_321 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_337 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_9_347 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_36 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_43 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_9_66 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_98 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_0 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_1 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_10 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_12 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_13 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_14 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_16 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_17 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_18 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_2 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_20 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_22 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_24 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_25 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_28 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_30 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_31 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_32 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_33 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_34 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_36 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_37 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_38 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_4 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_40 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_42 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_43 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_44 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_45 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_46 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_47 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_48 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_49 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_5 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_50 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_52 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_56 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_58 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_59 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_6 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_60 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_61 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_62 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_63 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_64 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_66 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_67 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_68 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_70 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_71 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_72 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_73 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_74 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_75 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_76 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_8 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_100 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_101 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_102 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_103 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_104 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_105 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_106 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_107 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_108 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_109 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_110 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_111 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_112 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_113 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_114 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_115 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_116 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_117 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_118 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_119 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_120 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_121 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_122 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_123 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_124 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_125 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_126 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_127 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_128 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_129 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_130 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_131 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_132 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_133 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_134 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_135 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_136 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_137 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_138 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_139 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_140 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_141 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_142 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_143 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_144 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_145 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_146 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_147 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_148 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_149 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_150 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_151 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_152 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_153 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_154 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_155 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_156 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_157 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_158 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_159 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_160 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_161 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_162 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_163 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_164 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_165 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_166 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_167 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_168 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_169 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_170 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_171 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_172 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_173 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_174 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_175 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_176 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_177 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_178 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_179 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_180 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_181 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_182 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_183 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_184 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_185 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_186 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_187 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_188 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_189 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_190 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_191 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_192 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_193 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_194 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_195 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_196 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_197 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_198 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_199 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_200 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_201 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_202 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_203 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_78 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_79 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_80 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_81 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_82 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_83 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_84 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_85 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_86 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_87 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_88 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_89 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_90 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_91 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_92 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_93 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_94 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_95 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_96 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_97 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_98 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_99 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__or3_1 _0469_ (.A(\u_driver.i_data[0] ),
    .B(\u_driver.i_data[3] ),
    .C(\u_driver.i_data[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0088_));
 sky130_fd_sc_hd__inv_2 _0470_ (.A(_0088_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0089_));
 sky130_fd_sc_hd__and3_1 _0471_ (.A(\u_driver.i_data[1] ),
    .B(\u_driver.i_valid ),
    .C(_0089_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0090_));
 sky130_fd_sc_hd__buf_1 _0472_ (.A(_0090_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\u_driver.dl_en ));
 sky130_fd_sc_hd__buf_2 _0473_ (.A(\u_tx.sm_uart_q[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0091_));
 sky130_fd_sc_hd__buf_2 _0474_ (.A(\u_tx.sm_uart_q[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0092_));
 sky130_fd_sc_hd__or3b_1 _0475_ (.A(\u_tx.sm_uart_q[3] ),
    .B(\u_tx.sm_uart_q[2] ),
    .C_N(\u_tx.sm_uart_q[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0093_));
 sky130_fd_sc_hd__a31o_1 _0476_ (.A1(_0091_),
    .A2(_0092_),
    .A3(\u_driver.data_edge[39] ),
    .B1(\u_tx.sm_uart_q[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0094_));
 sky130_fd_sc_hd__inv_2 _0477_ (.A(_0092_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0095_));
 sky130_fd_sc_hd__and3b_1 _0478_ (.A_N(_0091_),
    .B(_0092_),
    .C(\u_driver.data_edge[37] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0096_));
 sky130_fd_sc_hd__a31o_1 _0479_ (.A1(_0091_),
    .A2(_0095_),
    .A3(\u_driver.data_edge[38] ),
    .B1(_0096_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0097_));
 sky130_fd_sc_hd__and3b_1 _0480_ (.A_N(_0091_),
    .B(_0092_),
    .C(\u_driver.data_q[36] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0098_));
 sky130_fd_sc_hd__or3b_1 _0481_ (.A(_0091_),
    .B(_0092_),
    .C_N(\u_driver.data_in[39] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0099_));
 sky130_fd_sc_hd__nand2_1 _0482_ (.A(\u_tx.sm_uart_q[2] ),
    .B(_0099_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0100_));
 sky130_fd_sc_hd__a311o_1 _0483_ (.A1(_0091_),
    .A2(_0092_),
    .A3(\u_driver.data_q[38] ),
    .B1(_0098_),
    .C1(_0100_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0101_));
 sky130_fd_sc_hd__a31o_1 _0484_ (.A1(_0091_),
    .A2(_0095_),
    .A3(\u_driver.data_q[37] ),
    .B1(_0101_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0102_));
 sky130_fd_sc_hd__o21a_1 _0485_ (.A1(_0094_),
    .A2(_0097_),
    .B1(_0102_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0103_));
 sky130_fd_sc_hd__or3b_1 _0486_ (.A(\u_tx.sm_uart_q[4] ),
    .B(_0103_),
    .C_N(\u_tx.sm_uart_q[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0104_));
 sky130_fd_sc_hd__o41a_1 _0487_ (.A1(_0091_),
    .A2(_0092_),
    .A3(\u_driver.data_q[39] ),
    .A4(_0093_),
    .B1(_0104_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\u_tx.o_tx ));
 sky130_fd_sc_hd__or4b_1 _0488_ (.A(\u_rx.timer_q[1] ),
    .B(\u_rx.timer_q[0] ),
    .C(\u_rx.timer_q[2] ),
    .D_N(\u_rx.timer_q[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0105_));
 sky130_fd_sc_hd__or3_1 _0489_ (.A(\u_rx.timer_q[7] ),
    .B(\u_rx.timer_q[8] ),
    .C(_0105_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0106_));
 sky130_fd_sc_hd__inv_2 _0490_ (.A(\u_rx.timer_q[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0107_));
 sky130_fd_sc_hd__or4bb_1 _0491_ (.A(\u_rx.timer_q[5] ),
    .B(\u_rx.timer_q[9] ),
    .C_N(\u_rx.timer_q[6] ),
    .D_N(\u_rx.timer_q[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0108_));
 sky130_fd_sc_hd__or4b_1 _0492_ (.A(\u_rx.timer_q[11] ),
    .B(_0107_),
    .C(_0108_),
    .D_N(\u_rx.timer_q[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0109_));
 sky130_fd_sc_hd__inv_2 _0493_ (.A(\u_rx.sm_uart_q[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0110_));
 sky130_fd_sc_hd__or4b_1 _0494_ (.A(\u_rx.sm_uart_q[2] ),
    .B(_0110_),
    .C(net94),
    .D_N(\u_rx.sm_uart_q[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0111_));
 sky130_fd_sc_hd__nor3_1 _0495_ (.A(_0106_),
    .B(_0109_),
    .C(_0111_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_rx.valid_d ));
 sky130_fd_sc_hd__nor3b_1 _0496_ (.A(\u_driver.i_data[3] ),
    .B(\u_driver.i_data[2] ),
    .C_N(\u_driver.i_data[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0112_));
 sky130_fd_sc_hd__and3_2 _0497_ (.A(\u_driver.i_data[1] ),
    .B(\u_driver.i_valid ),
    .C(_0112_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0113_));
 sky130_fd_sc_hd__inv_2 _0498_ (.A(_0113_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0114_));
 sky130_fd_sc_hd__inv_2 _0499_ (.A(net48),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0115_));
 sky130_fd_sc_hd__nor2_1 _0500_ (.A(\u_driver.edge_cnt_q[0] ),
    .B(\u_driver.edge_cnt_q[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0116_));
 sky130_fd_sc_hd__and2b_1 _0501_ (.A_N(\u_driver.edge_cnt_q[2] ),
    .B(_0116_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0117_));
 sky130_fd_sc_hd__nand2_1 _0502_ (.A(_0115_),
    .B(_0117_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0118_));
 sky130_fd_sc_hd__nor2_2 _0503_ (.A(_0113_),
    .B(_0118_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0119_));
 sky130_fd_sc_hd__a21oi_1 _0504_ (.A1(net45),
    .A2(_0114_),
    .B1(_0119_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0000_));
 sky130_fd_sc_hd__and2_1 _0505_ (.A(\u_driver.edge_cnt_q[0] ),
    .B(\u_driver.edge_cnt_q[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0120_));
 sky130_fd_sc_hd__or2_1 _0506_ (.A(_0113_),
    .B(_0118_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0121_));
 sky130_fd_sc_hd__o31a_1 _0507_ (.A1(_0113_),
    .A2(_0116_),
    .A3(_0120_),
    .B1(_0121_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0001_));
 sky130_fd_sc_hd__o21a_1 _0508_ (.A1(\u_driver.edge_cnt_q[0] ),
    .A2(\u_driver.edge_cnt_q[1] ),
    .B1(\u_driver.edge_cnt_q[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0122_));
 sky130_fd_sc_hd__a211o_1 _0509_ (.A1(net48),
    .A2(_0117_),
    .B1(_0122_),
    .C1(_0113_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0002_));
 sky130_fd_sc_hd__o21ai_1 _0510_ (.A1(_0115_),
    .A2(_0117_),
    .B1(_0114_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0003_));
 sky130_fd_sc_hd__inv_2 _0511_ (.A(\u_driver.i_data[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0123_));
 sky130_fd_sc_hd__or4_1 _0512_ (.A(\u_tx.sm_uart_q[1] ),
    .B(\u_tx.sm_uart_q[0] ),
    .C(\u_tx.sm_uart_q[3] ),
    .D(\u_tx.sm_uart_q[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0124_));
 sky130_fd_sc_hd__nor2_2 _0513_ (.A(\u_tx.sm_uart_q[4] ),
    .B(_0124_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0125_));
 sky130_fd_sc_hd__inv_2 _0514_ (.A(\u_tx.timer_q[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0126_));
 sky130_fd_sc_hd__or4b_1 _0515_ (.A(\u_tx.timer_q[1] ),
    .B(\u_tx.timer_q[0] ),
    .C(\u_tx.timer_q[2] ),
    .D_N(\u_tx.timer_q[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0127_));
 sky130_fd_sc_hd__or4bb_1 _0516_ (.A(\u_tx.timer_q[7] ),
    .B(\u_tx.timer_q[9] ),
    .C_N(\u_tx.timer_q[12] ),
    .D_N(\u_tx.timer_q[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0128_));
 sky130_fd_sc_hd__or4b_1 _0517_ (.A(\u_tx.timer_q[8] ),
    .B(_0128_),
    .C(\u_tx.timer_q[11] ),
    .D_N(\u_tx.timer_q[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0129_));
 sky130_fd_sc_hd__or4_1 _0518_ (.A(\u_tx.timer_q[5] ),
    .B(_0126_),
    .C(_0127_),
    .D(_0129_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0130_));
 sky130_fd_sc_hd__nor2_2 _0519_ (.A(_0125_),
    .B(_0130_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0131_));
 sky130_fd_sc_hd__a21o_1 _0520_ (.A1(\u_driver.o_valid ),
    .A2(_0125_),
    .B1(_0131_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0132_));
 sky130_fd_sc_hd__and4bb_1 _0521_ (.A_N(_0093_),
    .B_N(\u_tx.sm_uart_q[1] ),
    .C(_0092_),
    .D(_0132_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0133_));
 sky130_fd_sc_hd__inv_2 _0522_ (.A(_0133_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0134_));
 sky130_fd_sc_hd__a32o_1 _0523_ (.A1(_0123_),
    .A2(\u_driver.i_valid ),
    .A3(_0112_),
    .B1(_0134_),
    .B2(net46),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0004_));
 sky130_fd_sc_hd__or2_2 _0524_ (.A(\u_tx.sm_uart_q[4] ),
    .B(_0124_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0135_));
 sky130_fd_sc_hd__and2_1 _0525_ (.A(_0135_),
    .B(_0130_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0136_));
 sky130_fd_sc_hd__mux2_1 _0526_ (.A0(_0136_),
    .A1(_0125_),
    .S(\u_tx.timer_q[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0137_));
 sky130_fd_sc_hd__clkbuf_1 _0527_ (.A(_0137_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0005_));
 sky130_fd_sc_hd__and3_1 _0528_ (.A(\u_tx.timer_q[1] ),
    .B(\u_tx.timer_q[0] ),
    .C(_0135_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0138_));
 sky130_fd_sc_hd__a21oi_1 _0529_ (.A1(\u_tx.timer_q[0] ),
    .A2(_0135_),
    .B1(net57),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0139_));
 sky130_fd_sc_hd__nor2_1 _0530_ (.A(_0138_),
    .B(net58),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0006_));
 sky130_fd_sc_hd__xor2_1 _0531_ (.A(net51),
    .B(_0138_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0007_));
 sky130_fd_sc_hd__and4_1 _0532_ (.A(\u_tx.timer_q[1] ),
    .B(\u_tx.timer_q[0] ),
    .C(\u_tx.timer_q[2] ),
    .D(\u_tx.timer_q[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0140_));
 sky130_fd_sc_hd__a21oi_1 _0533_ (.A1(\u_tx.timer_q[2] ),
    .A2(_0138_),
    .B1(net83),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0141_));
 sky130_fd_sc_hd__a211oi_1 _0534_ (.A1(_0135_),
    .A2(_0140_),
    .B1(net84),
    .C1(_0131_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0008_));
 sky130_fd_sc_hd__a21oi_1 _0535_ (.A1(_0135_),
    .A2(_0140_),
    .B1(\u_tx.timer_q[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0142_));
 sky130_fd_sc_hd__and3_1 _0536_ (.A(\u_tx.timer_q[4] ),
    .B(_0135_),
    .C(_0140_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0143_));
 sky130_fd_sc_hd__nor3_1 _0537_ (.A(_0131_),
    .B(_0142_),
    .C(_0143_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0009_));
 sky130_fd_sc_hd__xor2_1 _0538_ (.A(net59),
    .B(_0143_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0010_));
 sky130_fd_sc_hd__a31o_1 _0539_ (.A1(\u_tx.timer_q[5] ),
    .A2(\u_tx.timer_q[4] ),
    .A3(_0140_),
    .B1(\u_tx.timer_q[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0144_));
 sky130_fd_sc_hd__nand4_1 _0540_ (.A(\u_tx.timer_q[5] ),
    .B(\u_tx.timer_q[4] ),
    .C(\u_tx.timer_q[6] ),
    .D(_0140_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0145_));
 sky130_fd_sc_hd__a32o_1 _0541_ (.A1(_0136_),
    .A2(_0144_),
    .A3(_0145_),
    .B1(_0125_),
    .B2(net63),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0011_));
 sky130_fd_sc_hd__nor2_1 _0542_ (.A(_0125_),
    .B(_0145_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0146_));
 sky130_fd_sc_hd__xor2_1 _0543_ (.A(net55),
    .B(_0146_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0012_));
 sky130_fd_sc_hd__a21oi_1 _0544_ (.A1(\u_tx.timer_q[7] ),
    .A2(_0146_),
    .B1(net61),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0147_));
 sky130_fd_sc_hd__and3_1 _0545_ (.A(\u_tx.timer_q[7] ),
    .B(\u_tx.timer_q[8] ),
    .C(_0146_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0148_));
 sky130_fd_sc_hd__nor2_1 _0546_ (.A(net62),
    .B(_0148_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0013_));
 sky130_fd_sc_hd__xor2_1 _0547_ (.A(net52),
    .B(_0148_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0014_));
 sky130_fd_sc_hd__a21oi_1 _0548_ (.A1(\u_tx.timer_q[9] ),
    .A2(_0148_),
    .B1(net80),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0149_));
 sky130_fd_sc_hd__and3_1 _0549_ (.A(\u_tx.timer_q[9] ),
    .B(\u_tx.timer_q[10] ),
    .C(_0148_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0150_));
 sky130_fd_sc_hd__nor3_1 _0550_ (.A(_0131_),
    .B(_0149_),
    .C(_0150_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0015_));
 sky130_fd_sc_hd__xor2_1 _0551_ (.A(net50),
    .B(_0150_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0016_));
 sky130_fd_sc_hd__a21oi_1 _0552_ (.A1(\u_tx.timer_q[11] ),
    .A2(_0150_),
    .B1(net89),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0151_));
 sky130_fd_sc_hd__and3_1 _0553_ (.A(net89),
    .B(\u_tx.timer_q[11] ),
    .C(_0150_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0152_));
 sky130_fd_sc_hd__nor3_1 _0554_ (.A(_0131_),
    .B(_0151_),
    .C(_0152_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0017_));
 sky130_fd_sc_hd__or3_2 _0555_ (.A(\u_rx.sm_uart_q[2] ),
    .B(\u_rx.sm_uart_q[3] ),
    .C(\u_rx.sm_uart_q[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0153_));
 sky130_fd_sc_hd__or4b_1 _0556_ (.A(\u_rx.timer_q[7] ),
    .B(\u_rx.timer_q[8] ),
    .C(\u_rx.timer_q[9] ),
    .D_N(\u_rx.timer_q[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0154_));
 sky130_fd_sc_hd__or4b_1 _0557_ (.A(\u_rx.timer_q[11] ),
    .B(_0107_),
    .C(_0154_),
    .D_N(\u_rx.timer_q[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0155_));
 sky130_fd_sc_hd__or4bb_1 _0558_ (.A(\u_rx.timer_q[2] ),
    .B(\u_rx.timer_q[5] ),
    .C_N(\u_rx.timer_q[4] ),
    .D_N(\u_rx.timer_q[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0156_));
 sky130_fd_sc_hd__nor4_2 _0559_ (.A(\u_rx.timer_q[1] ),
    .B(\u_rx.timer_q[0] ),
    .C(_0155_),
    .D(_0156_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0157_));
 sky130_fd_sc_hd__nand2_4 _0560_ (.A(_0153_),
    .B(_0157_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0158_));
 sky130_fd_sc_hd__or4b_1 _0561_ (.A(\u_rx.sm_uart_q[1] ),
    .B(\u_rx.timer_q[1] ),
    .C(\u_rx.timer_q[0] ),
    .D_N(\u_rx.sm_uart_q[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0159_));
 sky130_fd_sc_hd__inv_2 _0562_ (.A(\u_rx.timer_q[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0160_));
 sky130_fd_sc_hd__nand2_1 _0563_ (.A(\u_rx.timer_q[3] ),
    .B(\u_rx.timer_q[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0161_));
 sky130_fd_sc_hd__or4b_1 _0564_ (.A(\u_rx.timer_q[7] ),
    .B(\u_rx.timer_q[6] ),
    .C(\u_rx.timer_q[8] ),
    .D_N(\u_rx.timer_q[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0162_));
 sky130_fd_sc_hd__or4b_1 _0565_ (.A(\u_rx.timer_q[10] ),
    .B(\u_rx.timer_q[12] ),
    .C(_0162_),
    .D_N(\u_rx.timer_q[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0163_));
 sky130_fd_sc_hd__or4_1 _0566_ (.A(\u_rx.timer_q[4] ),
    .B(_0160_),
    .C(_0161_),
    .D(_0163_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0164_));
 sky130_fd_sc_hd__nor4_1 _0567_ (.A(\u_rx.sm_uart_q[2] ),
    .B(\u_rx.sm_uart_q[3] ),
    .C(_0159_),
    .D(_0164_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0165_));
 sky130_fd_sc_hd__inv_2 _0568_ (.A(_0165_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0166_));
 sky130_fd_sc_hd__nand2_1 _0569_ (.A(_0158_),
    .B(_0166_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0167_));
 sky130_fd_sc_hd__o211a_1 _0570_ (.A1(\u_rx.sm_uart_q[0] ),
    .A2(_0153_),
    .B1(_0158_),
    .C1(_0166_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0168_));
 sky130_fd_sc_hd__inv_2 _0571_ (.A(net2),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0169_));
 sky130_fd_sc_hd__a211oi_2 _0572_ (.A1(\u_rx.p1_rx ),
    .A2(_0169_),
    .B1(\u_rx.sm_uart_q[0] ),
    .C1(_0153_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0170_));
 sky130_fd_sc_hd__clkbuf_4 _0573_ (.A(_0170_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0171_));
 sky130_fd_sc_hd__o21ba_1 _0574_ (.A1(_0168_),
    .A2(_0171_),
    .B1_N(\u_rx.sm_uart_q[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0172_));
 sky130_fd_sc_hd__a21oi_1 _0575_ (.A1(net66),
    .A2(_0167_),
    .B1(_0172_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0018_));
 sky130_fd_sc_hd__o211a_1 _0576_ (.A1(\u_rx.sm_uart_q[2] ),
    .A2(_0110_),
    .B1(\u_rx.sm_uart_q[0] ),
    .C1(_0167_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0173_));
 sky130_fd_sc_hd__and3_1 _0577_ (.A(\u_rx.sm_uart_q[1] ),
    .B(\u_rx.sm_uart_q[0] ),
    .C(_0167_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0174_));
 sky130_fd_sc_hd__o21ba_1 _0578_ (.A1(net67),
    .A2(_0173_),
    .B1_N(_0174_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0019_));
 sky130_fd_sc_hd__xor2_1 _0579_ (.A(net60),
    .B(_0174_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0020_));
 sky130_fd_sc_hd__a21oi_1 _0580_ (.A1(\u_rx.sm_uart_q[2] ),
    .A2(_0174_),
    .B1(\u_rx.sm_uart_q[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0175_));
 sky130_fd_sc_hd__and3_1 _0581_ (.A(\u_rx.sm_uart_q[2] ),
    .B(\u_rx.sm_uart_q[3] ),
    .C(_0174_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0176_));
 sky130_fd_sc_hd__or2_1 _0582_ (.A(_0175_),
    .B(_0176_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0177_));
 sky130_fd_sc_hd__and2b_1 _0583_ (.A_N(_0111_),
    .B(_0157_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0178_));
 sky130_fd_sc_hd__nor2_1 _0584_ (.A(_0177_),
    .B(_0178_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0021_));
 sky130_fd_sc_hd__mux2_1 _0585_ (.A0(\u_driver.i_data[1] ),
    .A1(net92),
    .S(_0158_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0179_));
 sky130_fd_sc_hd__clkbuf_1 _0586_ (.A(_0179_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0022_));
 sky130_fd_sc_hd__mux2_1 _0587_ (.A0(\u_driver.i_data[2] ),
    .A1(\u_driver.i_data[1] ),
    .S(_0158_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0180_));
 sky130_fd_sc_hd__clkbuf_1 _0588_ (.A(_0180_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0023_));
 sky130_fd_sc_hd__mux2_1 _0589_ (.A0(\u_driver.i_data[3] ),
    .A1(\u_driver.i_data[2] ),
    .S(_0158_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0181_));
 sky130_fd_sc_hd__clkbuf_1 _0590_ (.A(_0181_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0024_));
 sky130_fd_sc_hd__mux2_1 _0591_ (.A0(net78),
    .A1(\u_driver.i_data[3] ),
    .S(_0158_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0182_));
 sky130_fd_sc_hd__clkbuf_1 _0592_ (.A(_0182_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0025_));
 sky130_fd_sc_hd__mux2_1 _0593_ (.A0(\u_driver.data_in[1] ),
    .A1(\u_driver.data_in[0] ),
    .S(_0158_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0183_));
 sky130_fd_sc_hd__clkbuf_1 _0594_ (.A(_0183_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0026_));
 sky130_fd_sc_hd__mux2_1 _0595_ (.A0(\u_driver.data_in[2] ),
    .A1(\u_driver.data_in[1] ),
    .S(_0158_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0184_));
 sky130_fd_sc_hd__clkbuf_1 _0596_ (.A(_0184_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0027_));
 sky130_fd_sc_hd__mux2_1 _0597_ (.A0(\u_driver.data_in[3] ),
    .A1(\u_driver.data_in[2] ),
    .S(_0158_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0185_));
 sky130_fd_sc_hd__clkbuf_1 _0598_ (.A(_0185_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0028_));
 sky130_fd_sc_hd__mux2_1 _0599_ (.A0(net2),
    .A1(\u_driver.data_in[3] ),
    .S(_0158_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0186_));
 sky130_fd_sc_hd__clkbuf_1 _0600_ (.A(_0186_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0029_));
 sky130_fd_sc_hd__and2b_1 _0601_ (.A_N(\u_delay_line.data_4 ),
    .B(\u_delay_line.data_3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0187_));
 sky130_fd_sc_hd__or3b_1 _0602_ (.A(\u_delay_line.data_1 ),
    .B(_0187_),
    .C_N(\u_delay_line.data_0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0188_));
 sky130_fd_sc_hd__inv_2 _0603_ (.A(\u_delay_line.data_6 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0189_));
 sky130_fd_sc_hd__inv_2 _0604_ (.A(\u_delay_line.data_2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0190_));
 sky130_fd_sc_hd__o22a_1 _0605_ (.A1(\u_delay_line.data_7 ),
    .A2(_0189_),
    .B1(_0190_),
    .B2(\u_delay_line.data_3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0191_));
 sky130_fd_sc_hd__inv_2 _0606_ (.A(\u_delay_line.data_5 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0192_));
 sky130_fd_sc_hd__and2_1 _0607_ (.A(_0192_),
    .B(\u_delay_line.data_4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0193_));
 sky130_fd_sc_hd__inv_2 _0608_ (.A(_0193_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0194_));
 sky130_fd_sc_hd__inv_2 _0609_ (.A(\u_delay_line.data_8 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0195_));
 sky130_fd_sc_hd__inv_2 _0610_ (.A(\u_delay_line.data_9 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0196_));
 sky130_fd_sc_hd__nor2_1 _0611_ (.A(\u_delay_line.data_10 ),
    .B(_0196_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0197_));
 sky130_fd_sc_hd__a221o_1 _0612_ (.A1(_0195_),
    .A2(\u_delay_line.data_7 ),
    .B1(_0189_),
    .B2(\u_delay_line.data_5 ),
    .C1(_0197_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0198_));
 sky130_fd_sc_hd__a31o_1 _0613_ (.A1(_0188_),
    .A2(_0191_),
    .A3(_0194_),
    .B1(_0198_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0199_));
 sky130_fd_sc_hd__and2b_1 _0614_ (.A_N(\u_delay_line.data_11 ),
    .B(\u_delay_line.data_10 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0200_));
 sky130_fd_sc_hd__and2b_1 _0615_ (.A_N(\u_delay_line.data_13 ),
    .B(\u_delay_line.data_12 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0201_));
 sky130_fd_sc_hd__a211oi_1 _0616_ (.A1(\u_delay_line.data_8 ),
    .A2(_0196_),
    .B1(_0200_),
    .C1(_0201_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0202_));
 sky130_fd_sc_hd__and2b_1 _0617_ (.A_N(\u_delay_line.data_12 ),
    .B(\u_delay_line.data_11 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0203_));
 sky130_fd_sc_hd__and2b_1 _0618_ (.A_N(\u_delay_line.data_16 ),
    .B(\u_delay_line.data_15 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0204_));
 sky130_fd_sc_hd__and2b_1 _0619_ (.A_N(\u_delay_line.data_14 ),
    .B(\u_delay_line.data_13 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0205_));
 sky130_fd_sc_hd__or3_1 _0620_ (.A(_0203_),
    .B(_0204_),
    .C(_0205_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0206_));
 sky130_fd_sc_hd__a21oi_1 _0621_ (.A1(_0199_),
    .A2(_0202_),
    .B1(_0206_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0207_));
 sky130_fd_sc_hd__and2b_1 _0622_ (.A_N(\u_delay_line.data_19 ),
    .B(\u_delay_line.data_18 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0208_));
 sky130_fd_sc_hd__and2b_1 _0623_ (.A_N(\u_delay_line.data_15 ),
    .B(\u_delay_line.data_14 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0209_));
 sky130_fd_sc_hd__and2b_1 _0624_ (.A_N(\u_delay_line.data_17 ),
    .B(\u_delay_line.data_16 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0210_));
 sky130_fd_sc_hd__or4_1 _0625_ (.A(_0207_),
    .B(_0208_),
    .C(_0209_),
    .D(_0210_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0211_));
 sky130_fd_sc_hd__and2b_1 _0626_ (.A_N(\u_delay_line.data_18 ),
    .B(\u_delay_line.data_17 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0212_));
 sky130_fd_sc_hd__and2b_1 _0627_ (.A_N(\u_delay_line.data_22 ),
    .B(\u_delay_line.data_21 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0213_));
 sky130_fd_sc_hd__and2b_1 _0628_ (.A_N(\u_delay_line.data_20 ),
    .B(\u_delay_line.data_19 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0214_));
 sky130_fd_sc_hd__nor3_1 _0629_ (.A(_0212_),
    .B(_0213_),
    .C(_0214_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0215_));
 sky130_fd_sc_hd__and2b_1 _0630_ (.A_N(\u_delay_line.data_23 ),
    .B(\u_delay_line.data_22 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0216_));
 sky130_fd_sc_hd__and2b_1 _0631_ (.A_N(\u_delay_line.data_21 ),
    .B(\u_delay_line.data_20 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0217_));
 sky130_fd_sc_hd__and2b_1 _0632_ (.A_N(\u_delay_line.data_25 ),
    .B(\u_delay_line.data_24 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0218_));
 sky130_fd_sc_hd__or3_1 _0633_ (.A(_0216_),
    .B(_0217_),
    .C(_0218_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0219_));
 sky130_fd_sc_hd__a21o_1 _0634_ (.A1(_0211_),
    .A2(_0215_),
    .B1(_0219_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0220_));
 sky130_fd_sc_hd__inv_2 _0635_ (.A(\u_delay_line.data_26 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0221_));
 sky130_fd_sc_hd__nand2_1 _0636_ (.A(_0221_),
    .B(\u_delay_line.data_25 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0222_));
 sky130_fd_sc_hd__and2b_1 _0637_ (.A_N(\u_delay_line.data_28 ),
    .B(\u_delay_line.data_27 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0223_));
 sky130_fd_sc_hd__and2b_1 _0638_ (.A_N(\u_delay_line.data_24 ),
    .B(\u_delay_line.data_23 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0224_));
 sky130_fd_sc_hd__nor2_1 _0639_ (.A(_0223_),
    .B(_0224_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0225_));
 sky130_fd_sc_hd__inv_2 _0640_ (.A(\u_delay_line.data_31 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0226_));
 sky130_fd_sc_hd__inv_2 _0641_ (.A(\u_delay_line.data_29 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0227_));
 sky130_fd_sc_hd__and2_1 _0642_ (.A(\u_delay_line.data_28 ),
    .B(_0227_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0228_));
 sky130_fd_sc_hd__nor2_1 _0643_ (.A(_0221_),
    .B(\u_delay_line.data_27 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0229_));
 sky130_fd_sc_hd__a211o_1 _0644_ (.A1(\u_delay_line.data_30 ),
    .A2(_0226_),
    .B1(_0228_),
    .C1(_0229_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0230_));
 sky130_fd_sc_hd__a31o_1 _0645_ (.A1(_0220_),
    .A2(_0222_),
    .A3(_0225_),
    .B1(_0230_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0231_));
 sky130_fd_sc_hd__or2_1 _0646_ (.A(\u_driver.p1_capture ),
    .B(\u_driver.dl_en ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0232_));
 sky130_fd_sc_hd__buf_2 _0647_ (.A(_0232_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0233_));
 sky130_fd_sc_hd__nor2_2 _0648_ (.A(_0119_),
    .B(_0233_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0234_));
 sky130_fd_sc_hd__or2_1 _0649_ (.A(\u_delay_line.data_30 ),
    .B(_0227_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0235_));
 sky130_fd_sc_hd__a32o_1 _0650_ (.A1(_0231_),
    .A2(_0234_),
    .A3(_0235_),
    .B1(_0233_),
    .B2(\u_delay_line.data_0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0236_));
 sky130_fd_sc_hd__or3b_4 _0651_ (.A(_0088_),
    .B(\u_driver.i_data[1] ),
    .C_N(\u_driver.i_valid ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0237_));
 sky130_fd_sc_hd__mux2_1 _0652_ (.A0(\u_driver.data_in[0] ),
    .A1(_0236_),
    .S(_0237_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0238_));
 sky130_fd_sc_hd__and3_1 _0653_ (.A(_0123_),
    .B(\u_driver.i_valid ),
    .C(_0089_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0239_));
 sky130_fd_sc_hd__nor2_2 _0654_ (.A(\u_driver.p1_capture ),
    .B(\u_driver.dl_en ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0240_));
 sky130_fd_sc_hd__nand2_2 _0655_ (.A(_0119_),
    .B(_0240_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0241_));
 sky130_fd_sc_hd__a21o_1 _0656_ (.A1(\u_delay_line.valid_q ),
    .A2(_0241_),
    .B1(_0133_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0242_));
 sky130_fd_sc_hd__nor2_2 _0657_ (.A(_0239_),
    .B(_0242_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0243_));
 sky130_fd_sc_hd__clkbuf_4 _0658_ (.A(_0243_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0244_));
 sky130_fd_sc_hd__mux2_1 _0659_ (.A0(_0238_),
    .A1(\u_driver.data_dl[32] ),
    .S(_0244_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0245_));
 sky130_fd_sc_hd__clkbuf_1 _0660_ (.A(_0245_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0030_));
 sky130_fd_sc_hd__nand2_2 _0661_ (.A(_0121_),
    .B(_0240_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0246_));
 sky130_fd_sc_hd__clkbuf_4 _0662_ (.A(_0246_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0247_));
 sky130_fd_sc_hd__inv_2 _0663_ (.A(\u_delay_line.data_1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0248_));
 sky130_fd_sc_hd__mux2_1 _0664_ (.A0(\u_delay_line.data_3 ),
    .A1(_0248_),
    .S(_0190_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0249_));
 sky130_fd_sc_hd__mux2_1 _0665_ (.A0(\u_delay_line.data_7 ),
    .A1(_0192_),
    .S(_0189_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0250_));
 sky130_fd_sc_hd__o31a_1 _0666_ (.A1(_0187_),
    .A2(_0193_),
    .A3(_0249_),
    .B1(_0250_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0251_));
 sky130_fd_sc_hd__mux2_1 _0667_ (.A0(_0196_),
    .A1(\u_delay_line.data_7 ),
    .S(_0195_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0252_));
 sky130_fd_sc_hd__nor2_1 _0668_ (.A(_0197_),
    .B(_0200_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0253_));
 sky130_fd_sc_hd__o21a_1 _0669_ (.A1(_0251_),
    .A2(_0252_),
    .B1(_0253_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0254_));
 sky130_fd_sc_hd__nor2_1 _0670_ (.A(_0205_),
    .B(_0209_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0255_));
 sky130_fd_sc_hd__o31a_1 _0671_ (.A1(_0201_),
    .A2(_0203_),
    .A3(_0254_),
    .B1(_0255_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0256_));
 sky130_fd_sc_hd__or2_1 _0672_ (.A(_0204_),
    .B(_0210_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0257_));
 sky130_fd_sc_hd__nor2_1 _0673_ (.A(_0208_),
    .B(_0212_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0258_));
 sky130_fd_sc_hd__o21a_1 _0674_ (.A1(_0256_),
    .A2(_0257_),
    .B1(_0258_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0259_));
 sky130_fd_sc_hd__nor2_1 _0675_ (.A(_0213_),
    .B(_0216_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0260_));
 sky130_fd_sc_hd__o31a_1 _0676_ (.A1(_0214_),
    .A2(_0217_),
    .A3(_0259_),
    .B1(_0260_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0261_));
 sky130_fd_sc_hd__inv_2 _0677_ (.A(_0229_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0262_));
 sky130_fd_sc_hd__o311a_1 _0678_ (.A1(_0218_),
    .A2(_0224_),
    .A3(_0261_),
    .B1(_0262_),
    .C1(_0222_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0263_));
 sky130_fd_sc_hd__mux2_1 _0679_ (.A0(_0227_),
    .A1(\u_delay_line.data_31 ),
    .S(\u_delay_line.data_30 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0264_));
 sky130_fd_sc_hd__o31a_1 _0680_ (.A1(_0223_),
    .A2(_0228_),
    .A3(_0263_),
    .B1(_0264_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0265_));
 sky130_fd_sc_hd__nand2_1 _0681_ (.A(\u_delay_line.data_1 ),
    .B(_0233_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0266_));
 sky130_fd_sc_hd__o211a_1 _0682_ (.A1(_0247_),
    .A2(_0265_),
    .B1(_0266_),
    .C1(_0237_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0267_));
 sky130_fd_sc_hd__o21bai_1 _0683_ (.A1(\u_driver.data_in[1] ),
    .A2(_0237_),
    .B1_N(_0244_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0268_));
 sky130_fd_sc_hd__clkbuf_4 _0684_ (.A(_0243_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0269_));
 sky130_fd_sc_hd__a2bb2o_1 _0685_ (.A1_N(_0267_),
    .A2_N(_0268_),
    .B1(\u_driver.data_dl[33] ),
    .B2(_0269_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0031_));
 sky130_fd_sc_hd__or3b_1 _0686_ (.A(_0223_),
    .B(_0228_),
    .C_N(_0264_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0270_));
 sky130_fd_sc_hd__or4_1 _0687_ (.A(_0213_),
    .B(_0214_),
    .C(_0216_),
    .D(_0217_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0271_));
 sky130_fd_sc_hd__or4_1 _0688_ (.A(_0201_),
    .B(_0203_),
    .C(_0205_),
    .D(_0209_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0272_));
 sky130_fd_sc_hd__nor2_1 _0689_ (.A(_0187_),
    .B(_0193_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0273_));
 sky130_fd_sc_hd__or3_1 _0690_ (.A(_0197_),
    .B(_0200_),
    .C(_0252_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0274_));
 sky130_fd_sc_hd__a21oi_1 _0691_ (.A1(_0250_),
    .A2(_0273_),
    .B1(_0274_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0275_));
 sky130_fd_sc_hd__or3_1 _0692_ (.A(_0208_),
    .B(_0212_),
    .C(_0257_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0276_));
 sky130_fd_sc_hd__o21ba_1 _0693_ (.A1(_0272_),
    .A2(_0275_),
    .B1_N(_0276_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0277_));
 sky130_fd_sc_hd__a2111o_1 _0694_ (.A1(_0221_),
    .A2(\u_delay_line.data_25 ),
    .B1(_0218_),
    .C1(_0224_),
    .D1(_0229_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0278_));
 sky130_fd_sc_hd__o21ba_1 _0695_ (.A1(_0271_),
    .A2(_0277_),
    .B1_N(_0278_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0279_));
 sky130_fd_sc_hd__o21a_1 _0696_ (.A1(_0270_),
    .A2(_0279_),
    .B1(_0234_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0280_));
 sky130_fd_sc_hd__clkbuf_4 _0697_ (.A(_0239_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0281_));
 sky130_fd_sc_hd__a21o_1 _0698_ (.A1(\u_delay_line.data_2 ),
    .A2(_0233_),
    .B1(_0281_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0282_));
 sky130_fd_sc_hd__o22a_1 _0699_ (.A1(\u_driver.data_in[2] ),
    .A2(_0237_),
    .B1(_0280_),
    .B2(_0282_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0283_));
 sky130_fd_sc_hd__mux2_1 _0700_ (.A0(_0283_),
    .A1(\u_driver.data_dl[34] ),
    .S(_0244_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0284_));
 sky130_fd_sc_hd__clkbuf_1 _0701_ (.A(_0284_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0032_));
 sky130_fd_sc_hd__nor2_1 _0702_ (.A(_0270_),
    .B(_0278_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0285_));
 sky130_fd_sc_hd__nor2_1 _0703_ (.A(_0271_),
    .B(_0276_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0286_));
 sky130_fd_sc_hd__o21ai_1 _0704_ (.A1(_0272_),
    .A2(_0274_),
    .B1(_0286_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0287_));
 sky130_fd_sc_hd__a21oi_1 _0705_ (.A1(_0285_),
    .A2(_0287_),
    .B1(_0247_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0288_));
 sky130_fd_sc_hd__a21o_1 _0706_ (.A1(\u_delay_line.data_3 ),
    .A2(_0233_),
    .B1(_0281_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0289_));
 sky130_fd_sc_hd__o22a_1 _0707_ (.A1(\u_driver.data_in[3] ),
    .A2(_0237_),
    .B1(_0288_),
    .B2(_0289_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0290_));
 sky130_fd_sc_hd__mux2_1 _0708_ (.A0(_0290_),
    .A1(\u_driver.data_dl[35] ),
    .S(_0244_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0291_));
 sky130_fd_sc_hd__clkbuf_1 _0709_ (.A(_0291_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0033_));
 sky130_fd_sc_hd__a21oi_1 _0710_ (.A1(_0285_),
    .A2(_0286_),
    .B1(_0247_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0292_));
 sky130_fd_sc_hd__a21o_1 _0711_ (.A1(\u_delay_line.data_4 ),
    .A2(_0233_),
    .B1(_0281_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0293_));
 sky130_fd_sc_hd__o22a_1 _0712_ (.A1(\u_driver.data_dl[32] ),
    .A2(_0237_),
    .B1(_0292_),
    .B2(_0293_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0294_));
 sky130_fd_sc_hd__mux2_1 _0713_ (.A0(_0294_),
    .A1(\u_driver.data_dl[36] ),
    .S(_0244_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0295_));
 sky130_fd_sc_hd__clkbuf_1 _0714_ (.A(_0295_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0034_));
 sky130_fd_sc_hd__a22o_1 _0715_ (.A1(\u_delay_line.data_5 ),
    .A2(_0233_),
    .B1(_0234_),
    .B2(\u_driver.data_dl[32] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0296_));
 sky130_fd_sc_hd__and2_1 _0716_ (.A(_0237_),
    .B(_0242_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0297_));
 sky130_fd_sc_hd__buf_2 _0717_ (.A(_0297_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0298_));
 sky130_fd_sc_hd__clkbuf_4 _0718_ (.A(_0298_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0299_));
 sky130_fd_sc_hd__clkbuf_4 _0719_ (.A(_0239_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0300_));
 sky130_fd_sc_hd__and2_1 _0720_ (.A(\u_driver.data_dl[33] ),
    .B(_0300_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0301_));
 sky130_fd_sc_hd__a221o_1 _0721_ (.A1(net90),
    .A2(_0269_),
    .B1(_0296_),
    .B2(_0299_),
    .C1(_0301_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0035_));
 sky130_fd_sc_hd__a22o_1 _0722_ (.A1(\u_delay_line.data_6 ),
    .A2(_0233_),
    .B1(_0234_),
    .B2(\u_driver.data_dl[33] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0302_));
 sky130_fd_sc_hd__and2_1 _0723_ (.A(\u_driver.data_dl[34] ),
    .B(_0300_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0303_));
 sky130_fd_sc_hd__a221o_1 _0724_ (.A1(net88),
    .A2(_0269_),
    .B1(_0302_),
    .B2(_0299_),
    .C1(_0303_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0036_));
 sky130_fd_sc_hd__a22o_1 _0725_ (.A1(\u_delay_line.data_7 ),
    .A2(_0233_),
    .B1(_0234_),
    .B2(\u_driver.data_dl[34] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0304_));
 sky130_fd_sc_hd__and2_1 _0726_ (.A(\u_driver.data_dl[35] ),
    .B(_0300_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0305_));
 sky130_fd_sc_hd__a221o_1 _0727_ (.A1(net82),
    .A2(_0269_),
    .B1(_0304_),
    .B2(_0299_),
    .C1(_0305_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0037_));
 sky130_fd_sc_hd__clkbuf_4 _0728_ (.A(_0240_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0306_));
 sky130_fd_sc_hd__clkbuf_4 _0729_ (.A(_0246_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0307_));
 sky130_fd_sc_hd__buf_2 _0730_ (.A(_0241_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0308_));
 sky130_fd_sc_hd__o22a_1 _0731_ (.A1(\u_driver.data_dl[35] ),
    .A2(_0307_),
    .B1(_0308_),
    .B2(\u_driver.data_dl[32] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0309_));
 sky130_fd_sc_hd__o211a_1 _0732_ (.A1(\u_delay_line.data_8 ),
    .A2(_0306_),
    .B1(_0299_),
    .C1(_0309_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0310_));
 sky130_fd_sc_hd__a22o_1 _0733_ (.A1(\u_driver.data_dl[36] ),
    .A2(_0300_),
    .B1(_0244_),
    .B2(\u_driver.data_edge[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0311_));
 sky130_fd_sc_hd__or2_1 _0734_ (.A(_0310_),
    .B(_0311_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0312_));
 sky130_fd_sc_hd__clkbuf_1 _0735_ (.A(_0312_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0038_));
 sky130_fd_sc_hd__buf_2 _0736_ (.A(_0298_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0313_));
 sky130_fd_sc_hd__o22a_1 _0737_ (.A1(\u_driver.data_dl[36] ),
    .A2(_0307_),
    .B1(_0308_),
    .B2(\u_driver.data_dl[33] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0314_));
 sky130_fd_sc_hd__o211a_1 _0738_ (.A1(\u_delay_line.data_9 ),
    .A2(_0306_),
    .B1(_0313_),
    .C1(_0314_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0315_));
 sky130_fd_sc_hd__buf_2 _0739_ (.A(_0281_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0316_));
 sky130_fd_sc_hd__a22o_1 _0740_ (.A1(\u_driver.data_dl[37] ),
    .A2(_0316_),
    .B1(_0244_),
    .B2(\u_driver.data_edge[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0317_));
 sky130_fd_sc_hd__or2_1 _0741_ (.A(_0315_),
    .B(_0317_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0318_));
 sky130_fd_sc_hd__clkbuf_1 _0742_ (.A(_0318_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0039_));
 sky130_fd_sc_hd__o22a_1 _0743_ (.A1(\u_driver.data_dl[37] ),
    .A2(_0307_),
    .B1(_0308_),
    .B2(\u_driver.data_dl[34] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0319_));
 sky130_fd_sc_hd__o211a_1 _0744_ (.A1(\u_delay_line.data_10 ),
    .A2(_0306_),
    .B1(_0313_),
    .C1(_0319_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0320_));
 sky130_fd_sc_hd__a22o_1 _0745_ (.A1(\u_driver.data_dl[38] ),
    .A2(_0316_),
    .B1(_0244_),
    .B2(\u_driver.data_edge[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0321_));
 sky130_fd_sc_hd__or2_1 _0746_ (.A(_0320_),
    .B(_0321_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0322_));
 sky130_fd_sc_hd__clkbuf_1 _0747_ (.A(_0322_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0040_));
 sky130_fd_sc_hd__o22a_1 _0748_ (.A1(\u_driver.data_dl[38] ),
    .A2(_0307_),
    .B1(_0308_),
    .B2(\u_driver.data_dl[35] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0323_));
 sky130_fd_sc_hd__o211a_1 _0749_ (.A1(\u_delay_line.data_11 ),
    .A2(_0306_),
    .B1(_0313_),
    .C1(_0323_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0324_));
 sky130_fd_sc_hd__a22o_1 _0750_ (.A1(\u_driver.data_dl[39] ),
    .A2(_0316_),
    .B1(_0244_),
    .B2(\u_driver.data_edge[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0325_));
 sky130_fd_sc_hd__or2_1 _0751_ (.A(_0324_),
    .B(_0325_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0326_));
 sky130_fd_sc_hd__clkbuf_1 _0752_ (.A(_0326_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0041_));
 sky130_fd_sc_hd__o22a_1 _0753_ (.A1(\u_driver.data_dl[39] ),
    .A2(_0307_),
    .B1(_0308_),
    .B2(\u_driver.data_dl[36] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0327_));
 sky130_fd_sc_hd__o211a_1 _0754_ (.A1(\u_delay_line.data_12 ),
    .A2(_0306_),
    .B1(_0313_),
    .C1(_0327_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0328_));
 sky130_fd_sc_hd__a22o_1 _0755_ (.A1(\u_driver.data_edge[13] ),
    .A2(_0316_),
    .B1(_0244_),
    .B2(\u_driver.data_edge[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0329_));
 sky130_fd_sc_hd__or2_1 _0756_ (.A(_0328_),
    .B(_0329_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0330_));
 sky130_fd_sc_hd__clkbuf_1 _0757_ (.A(_0330_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0042_));
 sky130_fd_sc_hd__clkbuf_4 _0758_ (.A(_0240_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0331_));
 sky130_fd_sc_hd__o22a_1 _0759_ (.A1(\u_driver.data_edge[13] ),
    .A2(_0307_),
    .B1(_0308_),
    .B2(\u_driver.data_dl[37] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0332_));
 sky130_fd_sc_hd__o211a_1 _0760_ (.A1(\u_delay_line.data_13 ),
    .A2(_0331_),
    .B1(_0313_),
    .C1(_0332_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0333_));
 sky130_fd_sc_hd__clkbuf_4 _0761_ (.A(_0243_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0334_));
 sky130_fd_sc_hd__a22o_1 _0762_ (.A1(\u_driver.data_edge[14] ),
    .A2(_0316_),
    .B1(_0334_),
    .B2(\u_driver.data_edge[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0335_));
 sky130_fd_sc_hd__or2_1 _0763_ (.A(_0333_),
    .B(_0335_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0336_));
 sky130_fd_sc_hd__clkbuf_1 _0764_ (.A(_0336_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0043_));
 sky130_fd_sc_hd__o22a_1 _0765_ (.A1(\u_driver.data_edge[14] ),
    .A2(_0307_),
    .B1(_0308_),
    .B2(\u_driver.data_dl[38] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0337_));
 sky130_fd_sc_hd__o211a_1 _0766_ (.A1(\u_delay_line.data_14 ),
    .A2(_0331_),
    .B1(_0313_),
    .C1(_0337_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0338_));
 sky130_fd_sc_hd__a22o_1 _0767_ (.A1(\u_driver.data_edge[15] ),
    .A2(_0316_),
    .B1(_0334_),
    .B2(\u_driver.data_edge[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0339_));
 sky130_fd_sc_hd__or2_1 _0768_ (.A(_0338_),
    .B(_0339_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0340_));
 sky130_fd_sc_hd__clkbuf_1 _0769_ (.A(_0340_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0044_));
 sky130_fd_sc_hd__clkbuf_4 _0770_ (.A(_0241_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0341_));
 sky130_fd_sc_hd__clkbuf_4 _0771_ (.A(_0240_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0342_));
 sky130_fd_sc_hd__o22a_1 _0772_ (.A1(\u_delay_line.data_15 ),
    .A2(_0342_),
    .B1(_0247_),
    .B2(\u_driver.data_edge[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0343_));
 sky130_fd_sc_hd__o211a_1 _0773_ (.A1(\u_driver.data_dl[39] ),
    .A2(_0341_),
    .B1(_0313_),
    .C1(_0343_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0344_));
 sky130_fd_sc_hd__a22o_1 _0774_ (.A1(\u_driver.data_edge[16] ),
    .A2(_0316_),
    .B1(_0334_),
    .B2(\u_driver.data_edge[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0345_));
 sky130_fd_sc_hd__or2_1 _0775_ (.A(_0344_),
    .B(_0345_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0346_));
 sky130_fd_sc_hd__clkbuf_1 _0776_ (.A(_0346_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0045_));
 sky130_fd_sc_hd__clkbuf_4 _0777_ (.A(_0246_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0347_));
 sky130_fd_sc_hd__o22a_1 _0778_ (.A1(\u_driver.data_edge[16] ),
    .A2(_0347_),
    .B1(_0308_),
    .B2(\u_driver.data_edge[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0348_));
 sky130_fd_sc_hd__o211a_1 _0779_ (.A1(\u_delay_line.data_16 ),
    .A2(_0331_),
    .B1(_0313_),
    .C1(_0348_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0349_));
 sky130_fd_sc_hd__a22o_1 _0780_ (.A1(\u_driver.data_edge[17] ),
    .A2(_0316_),
    .B1(_0334_),
    .B2(\u_driver.data_edge[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0350_));
 sky130_fd_sc_hd__or2_1 _0781_ (.A(_0349_),
    .B(_0350_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0351_));
 sky130_fd_sc_hd__clkbuf_1 _0782_ (.A(_0351_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0046_));
 sky130_fd_sc_hd__o22a_1 _0783_ (.A1(\u_driver.data_edge[17] ),
    .A2(_0347_),
    .B1(_0308_),
    .B2(\u_driver.data_edge[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0352_));
 sky130_fd_sc_hd__o211a_1 _0784_ (.A1(\u_delay_line.data_17 ),
    .A2(_0331_),
    .B1(_0313_),
    .C1(_0352_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0353_));
 sky130_fd_sc_hd__a22o_1 _0785_ (.A1(\u_driver.data_edge[18] ),
    .A2(_0316_),
    .B1(_0334_),
    .B2(\u_driver.data_edge[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0354_));
 sky130_fd_sc_hd__or2_1 _0786_ (.A(_0353_),
    .B(_0354_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0355_));
 sky130_fd_sc_hd__clkbuf_1 _0787_ (.A(_0355_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0047_));
 sky130_fd_sc_hd__o22a_1 _0788_ (.A1(\u_driver.data_edge[18] ),
    .A2(_0247_),
    .B1(_0341_),
    .B2(\u_driver.data_edge[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0356_));
 sky130_fd_sc_hd__o211a_1 _0789_ (.A1(\u_delay_line.data_18 ),
    .A2(_0306_),
    .B1(_0299_),
    .C1(_0356_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0357_));
 sky130_fd_sc_hd__a221o_1 _0790_ (.A1(\u_driver.data_edge[19] ),
    .A2(_0300_),
    .B1(_0269_),
    .B2(net75),
    .C1(_0357_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0048_));
 sky130_fd_sc_hd__o22a_1 _0791_ (.A1(\u_delay_line.data_19 ),
    .A2(_0342_),
    .B1(_0307_),
    .B2(\u_driver.data_edge[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0358_));
 sky130_fd_sc_hd__o211a_1 _0792_ (.A1(\u_driver.data_edge[16] ),
    .A2(_0341_),
    .B1(_0313_),
    .C1(_0358_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0359_));
 sky130_fd_sc_hd__a22o_1 _0793_ (.A1(\u_driver.data_edge[20] ),
    .A2(_0316_),
    .B1(_0334_),
    .B2(\u_driver.data_edge[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0360_));
 sky130_fd_sc_hd__or2_1 _0794_ (.A(_0359_),
    .B(_0360_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0361_));
 sky130_fd_sc_hd__clkbuf_1 _0795_ (.A(_0361_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0049_));
 sky130_fd_sc_hd__o22a_1 _0796_ (.A1(\u_delay_line.data_20 ),
    .A2(_0342_),
    .B1(_0247_),
    .B2(\u_driver.data_edge[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0362_));
 sky130_fd_sc_hd__o211a_1 _0797_ (.A1(\u_driver.data_edge[17] ),
    .A2(_0341_),
    .B1(_0299_),
    .C1(_0362_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0363_));
 sky130_fd_sc_hd__a221o_1 _0798_ (.A1(\u_driver.data_edge[21] ),
    .A2(_0300_),
    .B1(_0269_),
    .B2(net77),
    .C1(_0363_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0050_));
 sky130_fd_sc_hd__clkbuf_4 _0799_ (.A(_0298_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0364_));
 sky130_fd_sc_hd__o22a_1 _0800_ (.A1(\u_driver.data_edge[21] ),
    .A2(_0347_),
    .B1(_0308_),
    .B2(\u_driver.data_edge[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0365_));
 sky130_fd_sc_hd__o211a_1 _0801_ (.A1(\u_delay_line.data_21 ),
    .A2(_0331_),
    .B1(_0364_),
    .C1(_0365_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0366_));
 sky130_fd_sc_hd__clkbuf_4 _0802_ (.A(_0281_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0367_));
 sky130_fd_sc_hd__a22o_1 _0803_ (.A1(\u_driver.data_edge[22] ),
    .A2(_0367_),
    .B1(_0334_),
    .B2(\u_driver.data_edge[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0368_));
 sky130_fd_sc_hd__or2_1 _0804_ (.A(_0366_),
    .B(_0368_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0369_));
 sky130_fd_sc_hd__clkbuf_1 _0805_ (.A(_0369_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0051_));
 sky130_fd_sc_hd__buf_2 _0806_ (.A(_0241_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0370_));
 sky130_fd_sc_hd__o22a_1 _0807_ (.A1(\u_driver.data_edge[22] ),
    .A2(_0347_),
    .B1(_0370_),
    .B2(\u_driver.data_edge[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0371_));
 sky130_fd_sc_hd__o211a_1 _0808_ (.A1(\u_delay_line.data_22 ),
    .A2(_0331_),
    .B1(_0364_),
    .C1(_0371_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0372_));
 sky130_fd_sc_hd__a22o_1 _0809_ (.A1(\u_driver.data_edge[23] ),
    .A2(_0367_),
    .B1(_0334_),
    .B2(\u_driver.data_edge[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0373_));
 sky130_fd_sc_hd__or2_1 _0810_ (.A(_0372_),
    .B(_0373_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0374_));
 sky130_fd_sc_hd__clkbuf_1 _0811_ (.A(_0374_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0052_));
 sky130_fd_sc_hd__o22a_1 _0812_ (.A1(\u_driver.data_edge[23] ),
    .A2(_0247_),
    .B1(_0341_),
    .B2(\u_driver.data_edge[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0375_));
 sky130_fd_sc_hd__o211a_1 _0813_ (.A1(\u_delay_line.data_23 ),
    .A2(_0306_),
    .B1(_0299_),
    .C1(_0375_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0376_));
 sky130_fd_sc_hd__a221o_1 _0814_ (.A1(net64),
    .A2(_0300_),
    .B1(_0269_),
    .B2(\u_driver.data_edge[28] ),
    .C1(_0376_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0053_));
 sky130_fd_sc_hd__o22a_1 _0815_ (.A1(\u_driver.data_edge[24] ),
    .A2(_0347_),
    .B1(_0370_),
    .B2(\u_driver.data_edge[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0377_));
 sky130_fd_sc_hd__o211a_1 _0816_ (.A1(\u_delay_line.data_24 ),
    .A2(_0331_),
    .B1(_0364_),
    .C1(_0377_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0378_));
 sky130_fd_sc_hd__a22o_1 _0817_ (.A1(\u_driver.data_edge[25] ),
    .A2(_0367_),
    .B1(_0334_),
    .B2(\u_driver.data_edge[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0379_));
 sky130_fd_sc_hd__or2_1 _0818_ (.A(_0378_),
    .B(_0379_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0380_));
 sky130_fd_sc_hd__clkbuf_1 _0819_ (.A(_0380_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0054_));
 sky130_fd_sc_hd__o22a_1 _0820_ (.A1(\u_driver.data_edge[25] ),
    .A2(_0347_),
    .B1(_0370_),
    .B2(\u_driver.data_edge[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0381_));
 sky130_fd_sc_hd__o211a_1 _0821_ (.A1(\u_delay_line.data_25 ),
    .A2(_0331_),
    .B1(_0364_),
    .C1(_0381_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0382_));
 sky130_fd_sc_hd__a22o_1 _0822_ (.A1(\u_driver.data_edge[26] ),
    .A2(_0367_),
    .B1(_0334_),
    .B2(\u_driver.data_edge[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0383_));
 sky130_fd_sc_hd__or2_1 _0823_ (.A(_0382_),
    .B(_0383_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0384_));
 sky130_fd_sc_hd__clkbuf_1 _0824_ (.A(_0384_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0055_));
 sky130_fd_sc_hd__o22a_1 _0825_ (.A1(\u_driver.data_edge[26] ),
    .A2(_0347_),
    .B1(_0370_),
    .B2(\u_driver.data_edge[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0385_));
 sky130_fd_sc_hd__o211a_1 _0826_ (.A1(\u_delay_line.data_26 ),
    .A2(_0331_),
    .B1(_0364_),
    .C1(_0385_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0386_));
 sky130_fd_sc_hd__buf_2 _0827_ (.A(_0243_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0387_));
 sky130_fd_sc_hd__a22o_1 _0828_ (.A1(\u_driver.data_edge[27] ),
    .A2(_0367_),
    .B1(_0387_),
    .B2(\u_driver.data_edge[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0388_));
 sky130_fd_sc_hd__or2_1 _0829_ (.A(_0386_),
    .B(_0388_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0389_));
 sky130_fd_sc_hd__clkbuf_1 _0830_ (.A(_0389_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0056_));
 sky130_fd_sc_hd__o22a_1 _0831_ (.A1(\u_driver.data_edge[27] ),
    .A2(_0347_),
    .B1(_0370_),
    .B2(\u_driver.data_edge[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0390_));
 sky130_fd_sc_hd__o211a_1 _0832_ (.A1(\u_delay_line.data_27 ),
    .A2(_0331_),
    .B1(_0364_),
    .C1(_0390_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0391_));
 sky130_fd_sc_hd__a22o_1 _0833_ (.A1(\u_driver.data_edge[28] ),
    .A2(_0367_),
    .B1(_0387_),
    .B2(\u_driver.data_edge[32] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0392_));
 sky130_fd_sc_hd__or2_1 _0834_ (.A(_0391_),
    .B(_0392_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0393_));
 sky130_fd_sc_hd__clkbuf_1 _0835_ (.A(_0393_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0057_));
 sky130_fd_sc_hd__o22a_1 _0836_ (.A1(\u_driver.data_edge[28] ),
    .A2(_0247_),
    .B1(_0341_),
    .B2(\u_driver.data_edge[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0394_));
 sky130_fd_sc_hd__o211a_1 _0837_ (.A1(\u_delay_line.data_28 ),
    .A2(_0306_),
    .B1(_0299_),
    .C1(_0394_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0395_));
 sky130_fd_sc_hd__a221o_1 _0838_ (.A1(net86),
    .A2(_0300_),
    .B1(_0269_),
    .B2(\u_driver.data_edge[33] ),
    .C1(_0395_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0058_));
 sky130_fd_sc_hd__o22a_1 _0839_ (.A1(\u_driver.data_edge[29] ),
    .A2(_0347_),
    .B1(_0370_),
    .B2(\u_driver.data_edge[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0396_));
 sky130_fd_sc_hd__o211a_1 _0840_ (.A1(\u_delay_line.data_29 ),
    .A2(_0342_),
    .B1(_0364_),
    .C1(_0396_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0397_));
 sky130_fd_sc_hd__a22o_1 _0841_ (.A1(\u_driver.data_edge[30] ),
    .A2(_0367_),
    .B1(_0387_),
    .B2(\u_driver.data_edge[34] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0398_));
 sky130_fd_sc_hd__or2_1 _0842_ (.A(_0397_),
    .B(_0398_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0399_));
 sky130_fd_sc_hd__clkbuf_1 _0843_ (.A(_0399_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0059_));
 sky130_fd_sc_hd__o22a_1 _0844_ (.A1(\u_driver.data_edge[30] ),
    .A2(_0247_),
    .B1(_0341_),
    .B2(\u_driver.data_edge[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0400_));
 sky130_fd_sc_hd__o211a_1 _0845_ (.A1(\u_delay_line.data_30 ),
    .A2(_0306_),
    .B1(_0299_),
    .C1(_0400_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0401_));
 sky130_fd_sc_hd__a221o_1 _0846_ (.A1(net79),
    .A2(_0300_),
    .B1(_0269_),
    .B2(net72),
    .C1(_0401_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0060_));
 sky130_fd_sc_hd__o22a_1 _0847_ (.A1(\u_delay_line.data_31 ),
    .A2(_0240_),
    .B1(_0307_),
    .B2(\u_driver.data_edge[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0402_));
 sky130_fd_sc_hd__o211a_1 _0848_ (.A1(\u_driver.data_edge[28] ),
    .A2(_0341_),
    .B1(_0364_),
    .C1(_0402_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0403_));
 sky130_fd_sc_hd__a22o_1 _0849_ (.A1(\u_driver.data_edge[32] ),
    .A2(_0367_),
    .B1(_0387_),
    .B2(\u_driver.data_edge[36] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0404_));
 sky130_fd_sc_hd__or2_1 _0850_ (.A(_0403_),
    .B(_0404_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0405_));
 sky130_fd_sc_hd__clkbuf_1 _0851_ (.A(_0405_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0061_));
 sky130_fd_sc_hd__o22a_1 _0852_ (.A1(\u_driver.data_edge[32] ),
    .A2(_0347_),
    .B1(_0370_),
    .B2(\u_driver.data_edge[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0406_));
 sky130_fd_sc_hd__o211a_1 _0853_ (.A1(\u_driver.data_dl[32] ),
    .A2(_0342_),
    .B1(_0364_),
    .C1(_0406_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0407_));
 sky130_fd_sc_hd__a22o_1 _0854_ (.A1(\u_driver.data_edge[33] ),
    .A2(_0367_),
    .B1(_0387_),
    .B2(\u_driver.data_edge[37] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0408_));
 sky130_fd_sc_hd__or2_1 _0855_ (.A(_0407_),
    .B(_0408_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0409_));
 sky130_fd_sc_hd__clkbuf_1 _0856_ (.A(_0409_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0062_));
 sky130_fd_sc_hd__o22a_1 _0857_ (.A1(\u_driver.data_edge[33] ),
    .A2(_0246_),
    .B1(_0370_),
    .B2(\u_driver.data_edge[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0410_));
 sky130_fd_sc_hd__o211a_1 _0858_ (.A1(\u_driver.data_dl[33] ),
    .A2(_0342_),
    .B1(_0364_),
    .C1(_0410_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0411_));
 sky130_fd_sc_hd__a22o_1 _0859_ (.A1(\u_driver.data_edge[34] ),
    .A2(_0367_),
    .B1(_0387_),
    .B2(\u_driver.data_edge[38] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0412_));
 sky130_fd_sc_hd__or2_1 _0860_ (.A(_0411_),
    .B(_0412_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0413_));
 sky130_fd_sc_hd__clkbuf_1 _0861_ (.A(_0413_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0063_));
 sky130_fd_sc_hd__o22a_1 _0862_ (.A1(\u_driver.data_edge[34] ),
    .A2(_0247_),
    .B1(_0341_),
    .B2(\u_driver.data_edge[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0414_));
 sky130_fd_sc_hd__o211a_1 _0863_ (.A1(\u_driver.data_dl[34] ),
    .A2(_0306_),
    .B1(_0299_),
    .C1(_0414_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0415_));
 sky130_fd_sc_hd__a221o_1 _0864_ (.A1(net72),
    .A2(_0300_),
    .B1(_0269_),
    .B2(\u_driver.data_edge[39] ),
    .C1(_0415_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0064_));
 sky130_fd_sc_hd__o22a_1 _0865_ (.A1(\u_driver.data_edge[35] ),
    .A2(_0246_),
    .B1(_0370_),
    .B2(\u_driver.data_edge[32] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0416_));
 sky130_fd_sc_hd__o211a_1 _0866_ (.A1(\u_driver.data_dl[35] ),
    .A2(_0342_),
    .B1(_0298_),
    .C1(_0416_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0417_));
 sky130_fd_sc_hd__a22o_1 _0867_ (.A1(\u_driver.data_edge[36] ),
    .A2(_0281_),
    .B1(_0387_),
    .B2(\u_driver.data_in[39] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0418_));
 sky130_fd_sc_hd__or2_1 _0868_ (.A(_0417_),
    .B(_0418_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0419_));
 sky130_fd_sc_hd__clkbuf_1 _0869_ (.A(_0419_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0065_));
 sky130_fd_sc_hd__o22a_1 _0870_ (.A1(\u_driver.data_dl[36] ),
    .A2(_0240_),
    .B1(_0307_),
    .B2(\u_driver.data_edge[36] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0420_));
 sky130_fd_sc_hd__o211a_1 _0871_ (.A1(\u_driver.data_edge[33] ),
    .A2(_0341_),
    .B1(_0298_),
    .C1(_0420_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0421_));
 sky130_fd_sc_hd__a22o_1 _0872_ (.A1(\u_driver.data_edge[37] ),
    .A2(_0281_),
    .B1(_0387_),
    .B2(\u_driver.data_q[36] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0422_));
 sky130_fd_sc_hd__or2_1 _0873_ (.A(_0421_),
    .B(_0422_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0423_));
 sky130_fd_sc_hd__clkbuf_1 _0874_ (.A(_0423_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0066_));
 sky130_fd_sc_hd__o22a_1 _0875_ (.A1(\u_driver.data_edge[37] ),
    .A2(_0246_),
    .B1(_0370_),
    .B2(\u_driver.data_edge[34] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0424_));
 sky130_fd_sc_hd__o211a_1 _0876_ (.A1(\u_driver.data_dl[37] ),
    .A2(_0342_),
    .B1(_0298_),
    .C1(_0424_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0425_));
 sky130_fd_sc_hd__a22o_1 _0877_ (.A1(\u_driver.data_edge[38] ),
    .A2(_0281_),
    .B1(_0387_),
    .B2(\u_driver.data_q[37] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0426_));
 sky130_fd_sc_hd__or2_1 _0878_ (.A(_0425_),
    .B(_0426_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0427_));
 sky130_fd_sc_hd__clkbuf_1 _0879_ (.A(_0427_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0067_));
 sky130_fd_sc_hd__o22a_1 _0880_ (.A1(\u_driver.data_edge[38] ),
    .A2(_0246_),
    .B1(_0241_),
    .B2(\u_driver.data_edge[35] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0428_));
 sky130_fd_sc_hd__o211a_1 _0881_ (.A1(\u_driver.data_dl[38] ),
    .A2(_0342_),
    .B1(_0298_),
    .C1(_0428_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0429_));
 sky130_fd_sc_hd__a22o_1 _0882_ (.A1(\u_driver.data_edge[39] ),
    .A2(_0281_),
    .B1(_0387_),
    .B2(\u_driver.data_q[38] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0430_));
 sky130_fd_sc_hd__or2_1 _0883_ (.A(_0429_),
    .B(_0430_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0431_));
 sky130_fd_sc_hd__clkbuf_1 _0884_ (.A(_0431_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0068_));
 sky130_fd_sc_hd__o22a_1 _0885_ (.A1(\u_driver.data_edge[39] ),
    .A2(_0246_),
    .B1(_0241_),
    .B2(\u_driver.data_edge[36] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0432_));
 sky130_fd_sc_hd__o211a_1 _0886_ (.A1(\u_driver.data_dl[39] ),
    .A2(_0342_),
    .B1(_0298_),
    .C1(_0432_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0433_));
 sky130_fd_sc_hd__a22o_1 _0887_ (.A1(\u_driver.data_in[39] ),
    .A2(_0281_),
    .B1(_0243_),
    .B2(\u_driver.data_q[39] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0434_));
 sky130_fd_sc_hd__or2_1 _0888_ (.A(_0433_),
    .B(_0434_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0435_));
 sky130_fd_sc_hd__clkbuf_1 _0889_ (.A(_0435_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0069_));
 sky130_fd_sc_hd__xnor2_1 _0890_ (.A(_0095_),
    .B(_0132_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0070_));
 sky130_fd_sc_hd__and3_1 _0891_ (.A(_0092_),
    .B(_0093_),
    .C(_0132_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0436_));
 sky130_fd_sc_hd__and3_1 _0892_ (.A(_0091_),
    .B(_0092_),
    .C(_0132_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0437_));
 sky130_fd_sc_hd__o21ba_1 _0893_ (.A1(_0091_),
    .A2(_0436_),
    .B1_N(_0437_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0071_));
 sky130_fd_sc_hd__nor2_1 _0894_ (.A(net93),
    .B(_0437_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0438_));
 sky130_fd_sc_hd__and2_1 _0895_ (.A(\u_tx.sm_uart_q[2] ),
    .B(_0437_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0439_));
 sky130_fd_sc_hd__nor2_1 _0896_ (.A(_0438_),
    .B(_0439_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0072_));
 sky130_fd_sc_hd__xor2_1 _0897_ (.A(net53),
    .B(_0439_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0073_));
 sky130_fd_sc_hd__a31o_1 _0898_ (.A1(\u_tx.sm_uart_q[3] ),
    .A2(\u_tx.sm_uart_q[2] ),
    .A3(_0437_),
    .B1(\u_tx.sm_uart_q[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0440_));
 sky130_fd_sc_hd__nand3_1 _0899_ (.A(\u_tx.sm_uart_q[4] ),
    .B(\u_tx.sm_uart_q[3] ),
    .C(_0439_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0441_));
 sky130_fd_sc_hd__and3_1 _0900_ (.A(_0134_),
    .B(_0440_),
    .C(_0441_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0442_));
 sky130_fd_sc_hd__clkbuf_1 _0901_ (.A(_0442_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0074_));
 sky130_fd_sc_hd__nor3_1 _0902_ (.A(_0157_),
    .B(_0165_),
    .C(_0170_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0443_));
 sky130_fd_sc_hd__clkbuf_4 _0903_ (.A(_0443_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0444_));
 sky130_fd_sc_hd__or2b_1 _0904_ (.A(_0170_),
    .B_N(\u_rx.timer_q[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0445_));
 sky130_fd_sc_hd__o21a_1 _0905_ (.A1(\u_rx.timer_q[0] ),
    .A2(_0444_),
    .B1(_0445_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0075_));
 sky130_fd_sc_hd__xnor2_1 _0906_ (.A(net85),
    .B(_0445_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0076_));
 sky130_fd_sc_hd__a21o_1 _0907_ (.A1(\u_rx.timer_q[1] ),
    .A2(\u_rx.timer_q[0] ),
    .B1(\u_rx.timer_q[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0446_));
 sky130_fd_sc_hd__nand3_1 _0908_ (.A(\u_rx.timer_q[1] ),
    .B(\u_rx.timer_q[0] ),
    .C(\u_rx.timer_q[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0447_));
 sky130_fd_sc_hd__a32o_1 _0909_ (.A1(_0444_),
    .A2(_0446_),
    .A3(_0447_),
    .B1(_0171_),
    .B2(net74),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0077_));
 sky130_fd_sc_hd__a31o_1 _0910_ (.A1(\u_rx.timer_q[1] ),
    .A2(\u_rx.timer_q[0] ),
    .A3(\u_rx.timer_q[2] ),
    .B1(\u_rx.timer_q[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0448_));
 sky130_fd_sc_hd__and4_1 _0911_ (.A(\u_rx.timer_q[1] ),
    .B(\u_rx.timer_q[0] ),
    .C(\u_rx.timer_q[3] ),
    .D(\u_rx.timer_q[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0449_));
 sky130_fd_sc_hd__inv_2 _0912_ (.A(_0449_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0450_));
 sky130_fd_sc_hd__a32o_1 _0913_ (.A1(_0444_),
    .A2(_0448_),
    .A3(_0450_),
    .B1(_0171_),
    .B2(net81),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0078_));
 sky130_fd_sc_hd__or2_1 _0914_ (.A(\u_rx.timer_q[4] ),
    .B(_0449_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0451_));
 sky130_fd_sc_hd__nand2_1 _0915_ (.A(\u_rx.timer_q[4] ),
    .B(_0449_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0452_));
 sky130_fd_sc_hd__a32o_1 _0916_ (.A1(_0444_),
    .A2(_0451_),
    .A3(_0452_),
    .B1(_0171_),
    .B2(net68),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0079_));
 sky130_fd_sc_hd__nand2_1 _0917_ (.A(_0160_),
    .B(_0452_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0453_));
 sky130_fd_sc_hd__nor2_1 _0918_ (.A(_0160_),
    .B(_0452_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0454_));
 sky130_fd_sc_hd__inv_2 _0919_ (.A(_0454_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0455_));
 sky130_fd_sc_hd__a32o_1 _0920_ (.A1(_0444_),
    .A2(_0453_),
    .A3(_0455_),
    .B1(_0171_),
    .B2(net71),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0080_));
 sky130_fd_sc_hd__and2_1 _0921_ (.A(\u_rx.timer_q[6] ),
    .B(_0454_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0456_));
 sky130_fd_sc_hd__o21ai_1 _0922_ (.A1(\u_rx.timer_q[6] ),
    .A2(_0454_),
    .B1(_0444_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0457_));
 sky130_fd_sc_hd__a2bb2o_1 _0923_ (.A1_N(_0456_),
    .A2_N(_0457_),
    .B1(net91),
    .B2(_0171_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0081_));
 sky130_fd_sc_hd__or2b_1 _0924_ (.A(_0170_),
    .B_N(_0456_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0458_));
 sky130_fd_sc_hd__xnor2_1 _0925_ (.A(net54),
    .B(_0458_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0082_));
 sky130_fd_sc_hd__and3b_1 _0926_ (.A_N(_0170_),
    .B(_0456_),
    .C(\u_rx.timer_q[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0459_));
 sky130_fd_sc_hd__xor2_1 _0927_ (.A(net56),
    .B(_0459_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0083_));
 sky130_fd_sc_hd__and4_2 _0928_ (.A(\u_rx.timer_q[7] ),
    .B(\u_rx.timer_q[8] ),
    .C(\u_rx.timer_q[9] ),
    .D(_0456_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0460_));
 sky130_fd_sc_hd__inv_2 _0929_ (.A(_0460_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0461_));
 sky130_fd_sc_hd__a31o_1 _0930_ (.A1(\u_rx.timer_q[7] ),
    .A2(\u_rx.timer_q[8] ),
    .A3(_0456_),
    .B1(\u_rx.timer_q[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0462_));
 sky130_fd_sc_hd__a32o_1 _0931_ (.A1(_0444_),
    .A2(_0461_),
    .A3(_0462_),
    .B1(_0171_),
    .B2(net70),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0084_));
 sky130_fd_sc_hd__nand2_1 _0932_ (.A(\u_rx.timer_q[10] ),
    .B(_0460_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0463_));
 sky130_fd_sc_hd__or2_1 _0933_ (.A(\u_rx.timer_q[10] ),
    .B(_0460_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0464_));
 sky130_fd_sc_hd__a32o_1 _0934_ (.A1(_0444_),
    .A2(_0463_),
    .A3(_0464_),
    .B1(_0171_),
    .B2(net69),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0085_));
 sky130_fd_sc_hd__and3_1 _0935_ (.A(\u_rx.timer_q[10] ),
    .B(\u_rx.timer_q[11] ),
    .C(_0460_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0465_));
 sky130_fd_sc_hd__and2b_1 _0936_ (.A_N(_0465_),
    .B(_0443_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0466_));
 sky130_fd_sc_hd__a31o_1 _0937_ (.A1(\u_rx.timer_q[10] ),
    .A2(_0444_),
    .A3(_0460_),
    .B1(\u_rx.timer_q[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0467_));
 sky130_fd_sc_hd__o21a_1 _0938_ (.A1(_0171_),
    .A2(_0466_),
    .B1(_0467_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0086_));
 sky130_fd_sc_hd__o21a_1 _0939_ (.A1(_0171_),
    .A2(_0466_),
    .B1(\u_rx.timer_q[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0468_));
 sky130_fd_sc_hd__a31o_1 _0940_ (.A1(_0107_),
    .A2(_0444_),
    .A3(_0465_),
    .B1(_0468_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0087_));
 sky130_fd_sc_hd__dfrtp_1 _0941_ (.CLK(clknet_4_11_0_clk),
    .D(_0000_),
    .RESET_B(net13),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\u_driver.edge_cnt_q[0] ));
 sky130_fd_sc_hd__dfrtp_1 _0942_ (.CLK(clknet_4_11_0_clk),
    .D(_0001_),
    .RESET_B(net13),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\u_driver.edge_cnt_q[1] ));
 sky130_fd_sc_hd__dfrtp_1 _0943_ (.CLK(clknet_4_11_0_clk),
    .D(net49),
    .RESET_B(net13),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\u_driver.edge_cnt_q[2] ));
 sky130_fd_sc_hd__dfrtp_1 _0944_ (.CLK(clknet_4_11_0_clk),
    .D(_0003_),
    .RESET_B(net13),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\u_driver.edge_cnt_q[3] ));
 sky130_fd_sc_hd__dfrtp_1 _0945_ (.CLK(clknet_4_14_0_clk),
    .D(net47),
    .RESET_B(net18),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\u_driver.o_valid ));
 sky130_fd_sc_hd__dfrtp_1 _0946_ (.CLK(clknet_4_7_0_clk),
    .D(net44),
    .RESET_B(net8),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\u_delay_line.start_q ));
 sky130_fd_sc_hd__dfrtp_1 _0947_ (.CLK(clknet_4_6_0_clk),
    .D(net43),
    .RESET_B(net8),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\u_delay_line.valid_q ));
 sky130_fd_sc_hd__dfrtp_1 _0948_ (.CLK(clknet_4_10_0_clk),
    .D(_0005_),
    .RESET_B(net12),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\u_tx.timer_q[0] ));
 sky130_fd_sc_hd__dfrtp_1 _0949_ (.CLK(clknet_4_11_0_clk),
    .D(_0006_),
    .RESET_B(net14),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\u_tx.timer_q[1] ));
 sky130_fd_sc_hd__dfrtp_1 _0950_ (.CLK(clknet_4_11_0_clk),
    .D(_0007_),
    .RESET_B(net14),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\u_tx.timer_q[2] ));
 sky130_fd_sc_hd__dfrtp_1 _0951_ (.CLK(clknet_4_10_0_clk),
    .D(_0008_),
    .RESET_B(net14),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\u_tx.timer_q[3] ));
 sky130_fd_sc_hd__dfrtp_2 _0952_ (.CLK(clknet_4_10_0_clk),
    .D(_0009_),
    .RESET_B(net12),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\u_tx.timer_q[4] ));
 sky130_fd_sc_hd__dfrtp_1 _0953_ (.CLK(clknet_4_10_0_clk),
    .D(_0010_),
    .RESET_B(net12),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\u_tx.timer_q[5] ));
 sky130_fd_sc_hd__dfrtp_1 _0954_ (.CLK(clknet_4_10_0_clk),
    .D(_0011_),
    .RESET_B(net12),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\u_tx.timer_q[6] ));
 sky130_fd_sc_hd__dfrtp_1 _0955_ (.CLK(clknet_4_10_0_clk),
    .D(_0012_),
    .RESET_B(net12),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\u_tx.timer_q[7] ));
 sky130_fd_sc_hd__dfrtp_1 _0956_ (.CLK(clknet_4_10_0_clk),
    .D(_0013_),
    .RESET_B(net12),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\u_tx.timer_q[8] ));
 sky130_fd_sc_hd__dfrtp_1 _0957_ (.CLK(clknet_4_10_0_clk),
    .D(_0014_),
    .RESET_B(net12),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\u_tx.timer_q[9] ));
 sky130_fd_sc_hd__dfrtp_1 _0958_ (.CLK(clknet_4_10_0_clk),
    .D(_0015_),
    .RESET_B(net14),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\u_tx.timer_q[10] ));
 sky130_fd_sc_hd__dfrtp_1 _0959_ (.CLK(clknet_4_10_0_clk),
    .D(_0016_),
    .RESET_B(net14),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\u_tx.timer_q[11] ));
 sky130_fd_sc_hd__dfrtp_1 _0960_ (.CLK(clknet_4_10_0_clk),
    .D(_0017_),
    .RESET_B(net14),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\u_tx.timer_q[12] ));
 sky130_fd_sc_hd__dfstp_1 _0961_ (.CLK(clknet_4_13_0_clk),
    .D(net2),
    .SET_B(net16),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\u_rx.p1_rx ));
 sky130_fd_sc_hd__dfrtp_4 _0962_ (.CLK(clknet_4_15_0_clk),
    .D(_0018_),
    .RESET_B(net18),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\u_rx.sm_uart_q[0] ));
 sky130_fd_sc_hd__dfrtp_1 _0963_ (.CLK(clknet_4_15_0_clk),
    .D(_0019_),
    .RESET_B(net19),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\u_rx.sm_uart_q[1] ));
 sky130_fd_sc_hd__dfrtp_2 _0964_ (.CLK(clknet_4_15_0_clk),
    .D(_0020_),
    .RESET_B(net19),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\u_rx.sm_uart_q[2] ));
 sky130_fd_sc_hd__dfrtp_1 _0965_ (.CLK(clknet_4_13_0_clk),
    .D(_0021_),
    .RESET_B(net16),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\u_rx.sm_uart_q[3] ));
 sky130_fd_sc_hd__dfrtp_1 _0966_ (.CLK(clknet_4_14_0_clk),
    .D(_0022_),
    .RESET_B(net16),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\u_driver.i_data[0] ));
 sky130_fd_sc_hd__dfrtp_2 _0967_ (.CLK(clknet_4_15_0_clk),
    .D(_0023_),
    .RESET_B(net19),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\u_driver.i_data[1] ));
 sky130_fd_sc_hd__dfrtp_1 _0968_ (.CLK(clknet_4_15_0_clk),
    .D(_0024_),
    .RESET_B(net19),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\u_driver.i_data[2] ));
 sky130_fd_sc_hd__dfrtp_1 _0969_ (.CLK(clknet_4_13_0_clk),
    .D(_0025_),
    .RESET_B(net17),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\u_driver.i_data[3] ));
 sky130_fd_sc_hd__dfrtp_1 _0970_ (.CLK(clknet_4_12_0_clk),
    .D(_0026_),
    .RESET_B(net16),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\u_driver.data_in[0] ));
 sky130_fd_sc_hd__dfrtp_1 _0971_ (.CLK(clknet_4_7_0_clk),
    .D(_0027_),
    .RESET_B(net16),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\u_driver.data_in[1] ));
 sky130_fd_sc_hd__dfrtp_1 _0972_ (.CLK(clknet_4_7_0_clk),
    .D(_0028_),
    .RESET_B(net8),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\u_driver.data_in[2] ));
 sky130_fd_sc_hd__dfrtp_1 _0973_ (.CLK(clknet_4_7_0_clk),
    .D(_0029_),
    .RESET_B(net8),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\u_driver.data_in[3] ));
 sky130_fd_sc_hd__dfrtp_1 _0974_ (.CLK(clknet_4_13_0_clk),
    .D(\u_rx.valid_d ),
    .RESET_B(net17),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\u_driver.i_valid ));
 sky130_fd_sc_hd__dfrtp_2 _0975_ (.CLK(clknet_4_12_0_clk),
    .D(_0030_),
    .RESET_B(net16),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\u_driver.data_dl[32] ));
 sky130_fd_sc_hd__dfrtp_2 _0976_ (.CLK(clknet_4_9_0_clk),
    .D(_0031_),
    .RESET_B(net11),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\u_driver.data_dl[33] ));
 sky130_fd_sc_hd__dfrtp_2 _0977_ (.CLK(clknet_4_3_0_clk),
    .D(_0032_),
    .RESET_B(net5),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\u_driver.data_dl[34] ));
 sky130_fd_sc_hd__dfrtp_2 _0978_ (.CLK(clknet_4_6_0_clk),
    .D(_0033_),
    .RESET_B(net8),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\u_driver.data_dl[35] ));
 sky130_fd_sc_hd__dfrtp_2 _0979_ (.CLK(clknet_4_6_0_clk),
    .D(_0034_),
    .RESET_B(net16),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\u_driver.data_dl[36] ));
 sky130_fd_sc_hd__dfrtp_2 _0980_ (.CLK(clknet_4_9_0_clk),
    .D(_0035_),
    .RESET_B(net11),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\u_driver.data_dl[37] ));
 sky130_fd_sc_hd__dfrtp_2 _0981_ (.CLK(clknet_4_12_0_clk),
    .D(_0036_),
    .RESET_B(net16),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\u_driver.data_dl[38] ));
 sky130_fd_sc_hd__dfrtp_2 _0982_ (.CLK(clknet_4_12_0_clk),
    .D(_0037_),
    .RESET_B(net16),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\u_driver.data_dl[39] ));
 sky130_fd_sc_hd__dfrtp_1 _0983_ (.CLK(clknet_4_6_0_clk),
    .D(_0038_),
    .RESET_B(net8),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\u_driver.data_edge[13] ));
 sky130_fd_sc_hd__dfrtp_1 _0984_ (.CLK(clknet_4_1_0_clk),
    .D(_0039_),
    .RESET_B(net5),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\u_driver.data_edge[14] ));
 sky130_fd_sc_hd__dfrtp_1 _0985_ (.CLK(clknet_4_4_0_clk),
    .D(_0040_),
    .RESET_B(net7),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\u_driver.data_edge[15] ));
 sky130_fd_sc_hd__dfrtp_1 _0986_ (.CLK(clknet_4_4_0_clk),
    .D(_0041_),
    .RESET_B(net8),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\u_driver.data_edge[16] ));
 sky130_fd_sc_hd__dfrtp_1 _0987_ (.CLK(clknet_4_6_0_clk),
    .D(_0042_),
    .RESET_B(net8),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\u_driver.data_edge[17] ));
 sky130_fd_sc_hd__dfrtp_1 _0988_ (.CLK(clknet_4_3_0_clk),
    .D(_0043_),
    .RESET_B(net5),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\u_driver.data_edge[18] ));
 sky130_fd_sc_hd__dfrtp_2 _0989_ (.CLK(clknet_4_1_0_clk),
    .D(_0044_),
    .RESET_B(net3),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\u_driver.data_edge[19] ));
 sky130_fd_sc_hd__dfrtp_1 _0990_ (.CLK(clknet_4_0_0_clk),
    .D(_0045_),
    .RESET_B(net3),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\u_driver.data_edge[20] ));
 sky130_fd_sc_hd__dfrtp_1 _0991_ (.CLK(clknet_4_0_0_clk),
    .D(_0046_),
    .RESET_B(net3),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\u_driver.data_edge[21] ));
 sky130_fd_sc_hd__dfrtp_1 _0992_ (.CLK(clknet_4_2_0_clk),
    .D(_0047_),
    .RESET_B(net5),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\u_driver.data_edge[22] ));
 sky130_fd_sc_hd__dfrtp_1 _0993_ (.CLK(clknet_4_3_0_clk),
    .D(net76),
    .RESET_B(net6),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\u_driver.data_edge[23] ));
 sky130_fd_sc_hd__dfrtp_1 _0994_ (.CLK(clknet_4_2_0_clk),
    .D(_0049_),
    .RESET_B(net5),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\u_driver.data_edge[24] ));
 sky130_fd_sc_hd__dfrtp_1 _0995_ (.CLK(clknet_4_3_0_clk),
    .D(_0050_),
    .RESET_B(net6),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\u_driver.data_edge[25] ));
 sky130_fd_sc_hd__dfrtp_1 _0996_ (.CLK(clknet_4_2_0_clk),
    .D(_0051_),
    .RESET_B(net5),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\u_driver.data_edge[26] ));
 sky130_fd_sc_hd__dfrtp_1 _0997_ (.CLK(clknet_4_8_0_clk),
    .D(_0052_),
    .RESET_B(net11),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\u_driver.data_edge[27] ));
 sky130_fd_sc_hd__dfrtp_1 _0998_ (.CLK(clknet_4_9_0_clk),
    .D(net65),
    .RESET_B(net11),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\u_driver.data_edge[28] ));
 sky130_fd_sc_hd__dfrtp_1 _0999_ (.CLK(clknet_4_8_0_clk),
    .D(_0054_),
    .RESET_B(net11),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\u_driver.data_edge[29] ));
 sky130_fd_sc_hd__dfrtp_1 _1000_ (.CLK(clknet_4_8_0_clk),
    .D(_0055_),
    .RESET_B(net11),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\u_driver.data_edge[30] ));
 sky130_fd_sc_hd__dfrtp_1 _1001_ (.CLK(clknet_4_8_0_clk),
    .D(_0056_),
    .RESET_B(net12),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\u_driver.data_edge[31] ));
 sky130_fd_sc_hd__dfrtp_1 _1002_ (.CLK(clknet_4_8_0_clk),
    .D(_0057_),
    .RESET_B(net12),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\u_driver.data_edge[32] ));
 sky130_fd_sc_hd__dfrtp_1 _1003_ (.CLK(clknet_4_9_0_clk),
    .D(net87),
    .RESET_B(net15),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\u_driver.data_edge[33] ));
 sky130_fd_sc_hd__dfrtp_1 _1004_ (.CLK(clknet_4_9_0_clk),
    .D(_0059_),
    .RESET_B(net13),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\u_driver.data_edge[34] ));
 sky130_fd_sc_hd__dfrtp_1 _1005_ (.CLK(clknet_4_9_0_clk),
    .D(_0060_),
    .RESET_B(net15),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\u_driver.data_edge[35] ));
 sky130_fd_sc_hd__dfrtp_1 _1006_ (.CLK(clknet_4_11_0_clk),
    .D(_0061_),
    .RESET_B(net13),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\u_driver.data_edge[36] ));
 sky130_fd_sc_hd__dfrtp_1 _1007_ (.CLK(clknet_4_9_0_clk),
    .D(_0062_),
    .RESET_B(net13),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\u_driver.data_edge[37] ));
 sky130_fd_sc_hd__dfrtp_1 _1008_ (.CLK(clknet_4_11_0_clk),
    .D(_0063_),
    .RESET_B(net13),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\u_driver.data_edge[38] ));
 sky130_fd_sc_hd__dfrtp_1 _1009_ (.CLK(clknet_4_12_0_clk),
    .D(net73),
    .RESET_B(net15),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\u_driver.data_edge[39] ));
 sky130_fd_sc_hd__dfrtp_1 _1010_ (.CLK(clknet_4_14_0_clk),
    .D(_0065_),
    .RESET_B(net18),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\u_driver.data_in[39] ));
 sky130_fd_sc_hd__dfrtp_1 _1011_ (.CLK(clknet_4_11_0_clk),
    .D(_0066_),
    .RESET_B(net13),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\u_driver.data_q[36] ));
 sky130_fd_sc_hd__dfrtp_1 _1012_ (.CLK(clknet_4_11_0_clk),
    .D(_0067_),
    .RESET_B(net13),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\u_driver.data_q[37] ));
 sky130_fd_sc_hd__dfrtp_1 _1013_ (.CLK(clknet_4_14_0_clk),
    .D(_0068_),
    .RESET_B(net18),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\u_driver.data_q[38] ));
 sky130_fd_sc_hd__dfrtp_1 _1014_ (.CLK(clknet_4_14_0_clk),
    .D(_0069_),
    .RESET_B(net18),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\u_driver.data_q[39] ));
 sky130_fd_sc_hd__dfrtp_1 _1015_ (.CLK(clknet_4_14_0_clk),
    .D(_0070_),
    .RESET_B(net18),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\u_tx.sm_uart_q[0] ));
 sky130_fd_sc_hd__dfrtp_1 _1016_ (.CLK(clknet_4_14_0_clk),
    .D(_0071_),
    .RESET_B(net18),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\u_tx.sm_uart_q[1] ));
 sky130_fd_sc_hd__dfrtp_2 _1017_ (.CLK(clknet_4_14_0_clk),
    .D(_0072_),
    .RESET_B(net18),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\u_tx.sm_uart_q[2] ));
 sky130_fd_sc_hd__dfrtp_1 _1018_ (.CLK(clknet_4_15_0_clk),
    .D(_0073_),
    .RESET_B(net18),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\u_tx.sm_uart_q[3] ));
 sky130_fd_sc_hd__dfrtp_2 _1019_ (.CLK(clknet_4_15_0_clk),
    .D(_0074_),
    .RESET_B(net18),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\u_tx.sm_uart_q[4] ));
 sky130_fd_sc_hd__dfrtp_4 _1020_ (.CLK(clknet_4_13_0_clk),
    .D(_0075_),
    .RESET_B(net17),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\u_rx.timer_q[0] ));
 sky130_fd_sc_hd__dfrtp_4 _1021_ (.CLK(clknet_4_13_0_clk),
    .D(_0076_),
    .RESET_B(net17),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\u_rx.timer_q[1] ));
 sky130_fd_sc_hd__dfrtp_2 _1022_ (.CLK(clknet_4_13_0_clk),
    .D(_0077_),
    .RESET_B(net17),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\u_rx.timer_q[2] ));
 sky130_fd_sc_hd__dfrtp_1 _1023_ (.CLK(clknet_4_7_0_clk),
    .D(_0078_),
    .RESET_B(net17),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\u_rx.timer_q[3] ));
 sky130_fd_sc_hd__dfrtp_1 _1024_ (.CLK(clknet_4_7_0_clk),
    .D(_0079_),
    .RESET_B(net8),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\u_rx.timer_q[4] ));
 sky130_fd_sc_hd__dfrtp_1 _1025_ (.CLK(clknet_4_7_0_clk),
    .D(_0080_),
    .RESET_B(net9),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\u_rx.timer_q[5] ));
 sky130_fd_sc_hd__dfrtp_1 _1026_ (.CLK(clknet_4_7_0_clk),
    .D(_0081_),
    .RESET_B(net9),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\u_rx.timer_q[6] ));
 sky130_fd_sc_hd__dfrtp_1 _1027_ (.CLK(clknet_4_13_0_clk),
    .D(_0082_),
    .RESET_B(net17),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\u_rx.timer_q[7] ));
 sky130_fd_sc_hd__dfrtp_1 _1028_ (.CLK(clknet_4_13_0_clk),
    .D(_0083_),
    .RESET_B(net17),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\u_rx.timer_q[8] ));
 sky130_fd_sc_hd__dfrtp_1 _1029_ (.CLK(clknet_4_7_0_clk),
    .D(_0084_),
    .RESET_B(net9),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\u_rx.timer_q[9] ));
 sky130_fd_sc_hd__dfrtp_2 _1030_ (.CLK(clknet_4_5_0_clk),
    .D(_0085_),
    .RESET_B(net9),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\u_rx.timer_q[10] ));
 sky130_fd_sc_hd__dfrtp_1 _1031_ (.CLK(clknet_4_5_0_clk),
    .D(_0086_),
    .RESET_B(net7),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\u_rx.timer_q[11] ));
 sky130_fd_sc_hd__dfrtp_1 _1032_ (.CLK(clknet_4_5_0_clk),
    .D(_0087_),
    .RESET_B(net10),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\u_rx.timer_q[12] ));
 sky130_fd_sc_hd__dfrtp_1 _1033_ (.CLK(clknet_4_12_0_clk),
    .D(\u_driver.dl_en ),
    .RESET_B(net16),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\u_driver.p1_capture ));
 sky130_fd_sc_hd__buf_2 _1057_ (.A(\u_delay_line.start_d ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\u_delay_line.u_bulk_0.dl_0 ));
 sky130_fd_sc_hd__buf_2 _1058_ (.A(net43),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\u_delay_line.valid_d ));
 sky130_fd_sc_hd__clkbuf_4 _1059_ (.A(\u_tx.o_tx ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[0]));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_4_0_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_4_10_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_4_11_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_4_12_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_4_13_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_4_14_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_4_15_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_4_1_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_4_2_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_4_3_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_4_4_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_4_5_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_4_6_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_4_7_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_4_8_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_4_9_0_clk));
 sky130_fd_sc_hd__clkbuf_2 fanout10 (.A(net1),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_4 fanout11 (.A(net15),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_4 fanout12 (.A(net14),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_4 fanout13 (.A(net14),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net13));
 sky130_fd_sc_hd__buf_2 fanout14 (.A(net15),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_2 fanout15 (.A(net1),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_4 fanout16 (.A(net19),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_4 fanout17 (.A(net19),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_4 fanout18 (.A(net19),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net18));
 sky130_fd_sc_hd__buf_2 fanout19 (.A(net1),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_4 fanout3 (.A(net6),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_2 fanout4 (.A(net6),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_4 fanout5 (.A(net6),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_2 fanout6 (.A(net1),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_4 fanout7 (.A(net10),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_4 fanout8 (.A(net10),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_2 fanout9 (.A(net10),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net9));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(\u_tx.timer_q[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net52));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(\u_tx.sm_uart_q[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net53));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(\u_rx.timer_q[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net54));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(\u_tx.timer_q[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net55));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(\u_rx.timer_q[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net56));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(\u_tx.timer_q[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net57));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(_0139_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net58));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(\u_tx.timer_q[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net59));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(\u_rx.sm_uart_q[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net60));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(\u_tx.timer_q[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net61));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(\u_delay_line.start_d ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net44));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(_0147_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net62));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(\u_tx.timer_q[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net63));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(\u_driver.data_edge[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net64));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(_0053_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net65));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(\u_rx.sm_uart_q[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net66));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(\u_rx.sm_uart_q[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net67));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(\u_rx.timer_q[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net68));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(\u_rx.timer_q[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net69));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(\u_rx.timer_q[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net70));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(\u_rx.timer_q[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net71));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(\u_driver.edge_cnt_q[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net45));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(\u_driver.data_edge[35] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net72));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(_0064_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net73));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(\u_rx.timer_q[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net74));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(\u_driver.data_edge[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net75));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(_0048_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net76));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(\u_driver.data_edge[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net77));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(\u_driver.data_in[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net78));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(\u_driver.data_edge[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net79));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(\u_tx.timer_q[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net80));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(\u_rx.timer_q[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net81));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(\u_driver.o_valid ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net46));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(\u_driver.data_dl[39] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net82));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(\u_tx.timer_q[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net83));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(_0141_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net84));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(\u_rx.timer_q[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net85));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(\u_driver.data_edge[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net86));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(_0058_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net87));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(\u_driver.data_dl[38] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net88));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(\u_tx.timer_q[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net89));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(\u_driver.data_dl[37] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net90));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(\u_rx.timer_q[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net91));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(_0004_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net47));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(\u_driver.i_data[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net92));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(\u_tx.sm_uart_q[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net93));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(\u_rx.sm_uart_q[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net94));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(\u_driver.edge_cnt_q[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net48));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(_0002_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net49));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(\u_tx.timer_q[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net50));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(\u_tx.timer_q[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net51));
 sky130_fd_sc_hd__buf_2 input1 (.A(rst_n),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_2 input2 (.A(ui_in[0]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 rebuffer1 (.A(\u_delay_line.start_q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net43));
 sky130_fd_sc_hd__conb_1 tt_um_ashleyjr_delay_line_20 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net20));
 sky130_fd_sc_hd__conb_1 tt_um_ashleyjr_delay_line_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net21));
 sky130_fd_sc_hd__conb_1 tt_um_ashleyjr_delay_line_22 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net22));
 sky130_fd_sc_hd__conb_1 tt_um_ashleyjr_delay_line_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net23));
 sky130_fd_sc_hd__conb_1 tt_um_ashleyjr_delay_line_24 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net24));
 sky130_fd_sc_hd__conb_1 tt_um_ashleyjr_delay_line_25 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net25));
 sky130_fd_sc_hd__conb_1 tt_um_ashleyjr_delay_line_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net26));
 sky130_fd_sc_hd__conb_1 tt_um_ashleyjr_delay_line_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net27));
 sky130_fd_sc_hd__conb_1 tt_um_ashleyjr_delay_line_28 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net28));
 sky130_fd_sc_hd__conb_1 tt_um_ashleyjr_delay_line_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net29));
 sky130_fd_sc_hd__conb_1 tt_um_ashleyjr_delay_line_30 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net30));
 sky130_fd_sc_hd__conb_1 tt_um_ashleyjr_delay_line_31 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net31));
 sky130_fd_sc_hd__conb_1 tt_um_ashleyjr_delay_line_32 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net32));
 sky130_fd_sc_hd__conb_1 tt_um_ashleyjr_delay_line_33 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net33));
 sky130_fd_sc_hd__conb_1 tt_um_ashleyjr_delay_line_34 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net34));
 sky130_fd_sc_hd__conb_1 tt_um_ashleyjr_delay_line_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net35));
 sky130_fd_sc_hd__conb_1 tt_um_ashleyjr_delay_line_36 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net36));
 sky130_fd_sc_hd__conb_1 tt_um_ashleyjr_delay_line_37 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net37));
 sky130_fd_sc_hd__conb_1 tt_um_ashleyjr_delay_line_38 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net38));
 sky130_fd_sc_hd__conb_1 tt_um_ashleyjr_delay_line_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net39));
 sky130_fd_sc_hd__conb_1 tt_um_ashleyjr_delay_line_40 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net40));
 sky130_fd_sc_hd__conb_1 tt_um_ashleyjr_delay_line_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net41));
 sky130_fd_sc_hd__conb_1 tt_um_ashleyjr_delay_line_42 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net42));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_0.u_inv_0  (.A(\u_delay_line.start_q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.start_d ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_0.u_inv_1  (.A(\u_delay_line.start_d ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_0.dl_1 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_0.u_inv_10  (.A(\u_delay_line.u_bulk_0.dl_9 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_0.dl_10 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_0.u_inv_11  (.A(\u_delay_line.u_bulk_0.dl_10 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_0.dl_11 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_0.u_inv_12  (.A(\u_delay_line.u_bulk_0.dl_11 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_0.dl_12 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_0.u_inv_13  (.A(\u_delay_line.u_bulk_0.dl_12 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_0.dl_13 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_0.u_inv_14  (.A(\u_delay_line.u_bulk_0.dl_13 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_0.dl_14 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_0.u_inv_15  (.A(\u_delay_line.u_bulk_0.dl_14 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.bulk_0 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_0.u_inv_2  (.A(\u_delay_line.u_bulk_0.dl_1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_0.dl_2 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_0.u_inv_3  (.A(\u_delay_line.u_bulk_0.dl_2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_0.dl_3 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_0.u_inv_4  (.A(\u_delay_line.u_bulk_0.dl_3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_0.dl_4 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_0.u_inv_5  (.A(\u_delay_line.u_bulk_0.dl_4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_0.dl_5 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_0.u_inv_6  (.A(\u_delay_line.u_bulk_0.dl_5 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_0.dl_6 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_0.u_inv_7  (.A(\u_delay_line.u_bulk_0.dl_6 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_0.dl_7 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_0.u_inv_8  (.A(\u_delay_line.u_bulk_0.dl_7 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_0.dl_8 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_0.u_inv_9  (.A(\u_delay_line.u_bulk_0.dl_8 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_0.dl_9 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_1.u_inv_0  (.A(\u_delay_line.bulk_0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_1.dl_0 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_1.u_inv_1  (.A(\u_delay_line.u_bulk_1.dl_0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_1.dl_1 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_1.u_inv_10  (.A(\u_delay_line.u_bulk_1.dl_9 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_1.dl_10 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_1.u_inv_11  (.A(\u_delay_line.u_bulk_1.dl_10 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_1.dl_11 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_1.u_inv_12  (.A(\u_delay_line.u_bulk_1.dl_11 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_1.dl_12 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_1.u_inv_13  (.A(\u_delay_line.u_bulk_1.dl_12 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_1.dl_13 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_1.u_inv_14  (.A(\u_delay_line.u_bulk_1.dl_13 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_1.dl_14 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_1.u_inv_15  (.A(\u_delay_line.u_bulk_1.dl_14 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.bulk_1 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_1.u_inv_2  (.A(\u_delay_line.u_bulk_1.dl_1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_1.dl_2 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_1.u_inv_3  (.A(\u_delay_line.u_bulk_1.dl_2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_1.dl_3 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_1.u_inv_4  (.A(\u_delay_line.u_bulk_1.dl_3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_1.dl_4 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_1.u_inv_5  (.A(\u_delay_line.u_bulk_1.dl_4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_1.dl_5 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_1.u_inv_6  (.A(\u_delay_line.u_bulk_1.dl_5 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_1.dl_6 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_1.u_inv_7  (.A(\u_delay_line.u_bulk_1.dl_6 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_1.dl_7 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_1.u_inv_8  (.A(\u_delay_line.u_bulk_1.dl_7 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_1.dl_8 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_1.u_inv_9  (.A(\u_delay_line.u_bulk_1.dl_8 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_1.dl_9 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_10.u_inv_0  (.A(\u_delay_line.bulk_9 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_10.dl_0 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_10.u_inv_1  (.A(\u_delay_line.u_bulk_10.dl_0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_10.dl_1 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_10.u_inv_10  (.A(\u_delay_line.u_bulk_10.dl_9 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_10.dl_10 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_10.u_inv_11  (.A(\u_delay_line.u_bulk_10.dl_10 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_10.dl_11 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_10.u_inv_12  (.A(\u_delay_line.u_bulk_10.dl_11 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_10.dl_12 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_10.u_inv_13  (.A(\u_delay_line.u_bulk_10.dl_12 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_10.dl_13 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_10.u_inv_14  (.A(\u_delay_line.u_bulk_10.dl_13 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_10.dl_14 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_10.u_inv_15  (.A(\u_delay_line.u_bulk_10.dl_14 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.bulk_10 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_10.u_inv_2  (.A(\u_delay_line.u_bulk_10.dl_1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_10.dl_2 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_10.u_inv_3  (.A(\u_delay_line.u_bulk_10.dl_2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_10.dl_3 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_10.u_inv_4  (.A(\u_delay_line.u_bulk_10.dl_3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_10.dl_4 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_10.u_inv_5  (.A(\u_delay_line.u_bulk_10.dl_4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_10.dl_5 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_10.u_inv_6  (.A(\u_delay_line.u_bulk_10.dl_5 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_10.dl_6 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_10.u_inv_7  (.A(\u_delay_line.u_bulk_10.dl_6 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_10.dl_7 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_10.u_inv_8  (.A(\u_delay_line.u_bulk_10.dl_7 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_10.dl_8 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_10.u_inv_9  (.A(\u_delay_line.u_bulk_10.dl_8 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_10.dl_9 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_11.u_inv_0  (.A(\u_delay_line.bulk_10 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_11.dl_0 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_11.u_inv_1  (.A(\u_delay_line.u_bulk_11.dl_0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_11.dl_1 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_11.u_inv_10  (.A(\u_delay_line.u_bulk_11.dl_9 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_11.dl_10 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_11.u_inv_11  (.A(\u_delay_line.u_bulk_11.dl_10 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_11.dl_11 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_11.u_inv_12  (.A(\u_delay_line.u_bulk_11.dl_11 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_11.dl_12 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_11.u_inv_13  (.A(\u_delay_line.u_bulk_11.dl_12 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_11.dl_13 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_11.u_inv_14  (.A(\u_delay_line.u_bulk_11.dl_13 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_11.dl_14 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_11.u_inv_15  (.A(\u_delay_line.u_bulk_11.dl_14 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.bulk_11 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_11.u_inv_2  (.A(\u_delay_line.u_bulk_11.dl_1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_11.dl_2 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_11.u_inv_3  (.A(\u_delay_line.u_bulk_11.dl_2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_11.dl_3 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_11.u_inv_4  (.A(\u_delay_line.u_bulk_11.dl_3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_11.dl_4 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_11.u_inv_5  (.A(\u_delay_line.u_bulk_11.dl_4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_11.dl_5 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_11.u_inv_6  (.A(\u_delay_line.u_bulk_11.dl_5 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_11.dl_6 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_11.u_inv_7  (.A(\u_delay_line.u_bulk_11.dl_6 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_11.dl_7 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_11.u_inv_8  (.A(\u_delay_line.u_bulk_11.dl_7 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_11.dl_8 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_11.u_inv_9  (.A(\u_delay_line.u_bulk_11.dl_8 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_11.dl_9 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_12.u_inv_0  (.A(\u_delay_line.bulk_11 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_12.dl_0 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_12.u_inv_1  (.A(\u_delay_line.u_bulk_12.dl_0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_12.dl_1 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_12.u_inv_10  (.A(\u_delay_line.u_bulk_12.dl_9 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_12.dl_10 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_12.u_inv_11  (.A(\u_delay_line.u_bulk_12.dl_10 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_12.dl_11 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_12.u_inv_12  (.A(\u_delay_line.u_bulk_12.dl_11 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_12.dl_12 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_12.u_inv_13  (.A(\u_delay_line.u_bulk_12.dl_12 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_12.dl_13 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_12.u_inv_14  (.A(\u_delay_line.u_bulk_12.dl_13 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_12.dl_14 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_12.u_inv_15  (.A(\u_delay_line.u_bulk_12.dl_14 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.bulk_12 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_12.u_inv_2  (.A(\u_delay_line.u_bulk_12.dl_1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_12.dl_2 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_12.u_inv_3  (.A(\u_delay_line.u_bulk_12.dl_2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_12.dl_3 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_12.u_inv_4  (.A(\u_delay_line.u_bulk_12.dl_3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_12.dl_4 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_12.u_inv_5  (.A(\u_delay_line.u_bulk_12.dl_4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_12.dl_5 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_12.u_inv_6  (.A(\u_delay_line.u_bulk_12.dl_5 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_12.dl_6 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_12.u_inv_7  (.A(\u_delay_line.u_bulk_12.dl_6 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_12.dl_7 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_12.u_inv_8  (.A(\u_delay_line.u_bulk_12.dl_7 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_12.dl_8 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_12.u_inv_9  (.A(\u_delay_line.u_bulk_12.dl_8 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_12.dl_9 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_13.u_inv_0  (.A(\u_delay_line.bulk_12 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_13.dl_0 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_13.u_inv_1  (.A(\u_delay_line.u_bulk_13.dl_0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_13.dl_1 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_13.u_inv_10  (.A(\u_delay_line.u_bulk_13.dl_9 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_13.dl_10 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_13.u_inv_11  (.A(\u_delay_line.u_bulk_13.dl_10 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_13.dl_11 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_13.u_inv_12  (.A(\u_delay_line.u_bulk_13.dl_11 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_13.dl_12 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_13.u_inv_13  (.A(\u_delay_line.u_bulk_13.dl_12 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_13.dl_13 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_13.u_inv_14  (.A(\u_delay_line.u_bulk_13.dl_13 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_13.dl_14 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_13.u_inv_15  (.A(\u_delay_line.u_bulk_13.dl_14 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.bulk_13 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_13.u_inv_2  (.A(\u_delay_line.u_bulk_13.dl_1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_13.dl_2 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_13.u_inv_3  (.A(\u_delay_line.u_bulk_13.dl_2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_13.dl_3 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_13.u_inv_4  (.A(\u_delay_line.u_bulk_13.dl_3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_13.dl_4 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_13.u_inv_5  (.A(\u_delay_line.u_bulk_13.dl_4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_13.dl_5 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_13.u_inv_6  (.A(\u_delay_line.u_bulk_13.dl_5 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_13.dl_6 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_13.u_inv_7  (.A(\u_delay_line.u_bulk_13.dl_6 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_13.dl_7 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_13.u_inv_8  (.A(\u_delay_line.u_bulk_13.dl_7 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_13.dl_8 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_13.u_inv_9  (.A(\u_delay_line.u_bulk_13.dl_8 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_13.dl_9 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_14.u_inv_0  (.A(\u_delay_line.bulk_13 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_14.dl_0 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_14.u_inv_1  (.A(\u_delay_line.u_bulk_14.dl_0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_14.dl_1 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_14.u_inv_10  (.A(\u_delay_line.u_bulk_14.dl_9 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_14.dl_10 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_14.u_inv_11  (.A(\u_delay_line.u_bulk_14.dl_10 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_14.dl_11 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_14.u_inv_12  (.A(\u_delay_line.u_bulk_14.dl_11 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_14.dl_12 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_14.u_inv_13  (.A(\u_delay_line.u_bulk_14.dl_12 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_14.dl_13 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_14.u_inv_14  (.A(\u_delay_line.u_bulk_14.dl_13 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_14.dl_14 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_14.u_inv_15  (.A(\u_delay_line.u_bulk_14.dl_14 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.bulk_14 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_14.u_inv_2  (.A(\u_delay_line.u_bulk_14.dl_1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_14.dl_2 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_14.u_inv_3  (.A(\u_delay_line.u_bulk_14.dl_2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_14.dl_3 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_14.u_inv_4  (.A(\u_delay_line.u_bulk_14.dl_3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_14.dl_4 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_14.u_inv_5  (.A(\u_delay_line.u_bulk_14.dl_4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_14.dl_5 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_14.u_inv_6  (.A(\u_delay_line.u_bulk_14.dl_5 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_14.dl_6 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_14.u_inv_7  (.A(\u_delay_line.u_bulk_14.dl_6 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_14.dl_7 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_14.u_inv_8  (.A(\u_delay_line.u_bulk_14.dl_7 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_14.dl_8 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_14.u_inv_9  (.A(\u_delay_line.u_bulk_14.dl_8 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_14.dl_9 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_15.u_inv_0  (.A(\u_delay_line.bulk_14 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_15.dl_0 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_15.u_inv_1  (.A(\u_delay_line.u_bulk_15.dl_0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_15.dl_1 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_15.u_inv_10  (.A(\u_delay_line.u_bulk_15.dl_9 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_15.dl_10 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_15.u_inv_11  (.A(\u_delay_line.u_bulk_15.dl_10 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_15.dl_11 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_15.u_inv_12  (.A(\u_delay_line.u_bulk_15.dl_11 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_15.dl_12 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_15.u_inv_13  (.A(\u_delay_line.u_bulk_15.dl_12 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_15.dl_13 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_15.u_inv_14  (.A(\u_delay_line.u_bulk_15.dl_13 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_15.dl_14 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_15.u_inv_15  (.A(\u_delay_line.u_bulk_15.dl_14 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.bulk_15 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_15.u_inv_2  (.A(\u_delay_line.u_bulk_15.dl_1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_15.dl_2 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_15.u_inv_3  (.A(\u_delay_line.u_bulk_15.dl_2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_15.dl_3 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_15.u_inv_4  (.A(\u_delay_line.u_bulk_15.dl_3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_15.dl_4 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_15.u_inv_5  (.A(\u_delay_line.u_bulk_15.dl_4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_15.dl_5 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_15.u_inv_6  (.A(\u_delay_line.u_bulk_15.dl_5 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_15.dl_6 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_15.u_inv_7  (.A(\u_delay_line.u_bulk_15.dl_6 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_15.dl_7 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_15.u_inv_8  (.A(\u_delay_line.u_bulk_15.dl_7 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_15.dl_8 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_15.u_inv_9  (.A(\u_delay_line.u_bulk_15.dl_8 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_15.dl_9 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_16.u_inv_0  (.A(\u_delay_line.bulk_15 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_16.dl_0 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_16.u_inv_1  (.A(\u_delay_line.u_bulk_16.dl_0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_16.dl_1 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_16.u_inv_10  (.A(\u_delay_line.u_bulk_16.dl_9 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_16.dl_10 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_16.u_inv_11  (.A(\u_delay_line.u_bulk_16.dl_10 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_16.dl_11 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_16.u_inv_12  (.A(\u_delay_line.u_bulk_16.dl_11 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_16.dl_12 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_16.u_inv_13  (.A(\u_delay_line.u_bulk_16.dl_12 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_16.dl_13 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_16.u_inv_14  (.A(\u_delay_line.u_bulk_16.dl_13 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_16.dl_14 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_16.u_inv_15  (.A(\u_delay_line.u_bulk_16.dl_14 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.bulk_16 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_16.u_inv_2  (.A(\u_delay_line.u_bulk_16.dl_1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_16.dl_2 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_16.u_inv_3  (.A(\u_delay_line.u_bulk_16.dl_2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_16.dl_3 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_16.u_inv_4  (.A(\u_delay_line.u_bulk_16.dl_3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_16.dl_4 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_16.u_inv_5  (.A(\u_delay_line.u_bulk_16.dl_4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_16.dl_5 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_16.u_inv_6  (.A(\u_delay_line.u_bulk_16.dl_5 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_16.dl_6 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_16.u_inv_7  (.A(\u_delay_line.u_bulk_16.dl_6 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_16.dl_7 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_16.u_inv_8  (.A(\u_delay_line.u_bulk_16.dl_7 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_16.dl_8 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_16.u_inv_9  (.A(\u_delay_line.u_bulk_16.dl_8 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_16.dl_9 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_17.u_inv_0  (.A(\u_delay_line.bulk_16 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_17.dl_0 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_17.u_inv_1  (.A(\u_delay_line.u_bulk_17.dl_0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_17.dl_1 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_17.u_inv_10  (.A(\u_delay_line.u_bulk_17.dl_9 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_17.dl_10 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_17.u_inv_11  (.A(\u_delay_line.u_bulk_17.dl_10 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_17.dl_11 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_17.u_inv_12  (.A(\u_delay_line.u_bulk_17.dl_11 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_17.dl_12 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_17.u_inv_13  (.A(\u_delay_line.u_bulk_17.dl_12 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_17.dl_13 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_17.u_inv_14  (.A(\u_delay_line.u_bulk_17.dl_13 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_17.dl_14 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_17.u_inv_15  (.A(\u_delay_line.u_bulk_17.dl_14 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.bulk_17 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_17.u_inv_2  (.A(\u_delay_line.u_bulk_17.dl_1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_17.dl_2 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_17.u_inv_3  (.A(\u_delay_line.u_bulk_17.dl_2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_17.dl_3 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_17.u_inv_4  (.A(\u_delay_line.u_bulk_17.dl_3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_17.dl_4 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_17.u_inv_5  (.A(\u_delay_line.u_bulk_17.dl_4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_17.dl_5 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_17.u_inv_6  (.A(\u_delay_line.u_bulk_17.dl_5 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_17.dl_6 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_17.u_inv_7  (.A(\u_delay_line.u_bulk_17.dl_6 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_17.dl_7 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_17.u_inv_8  (.A(\u_delay_line.u_bulk_17.dl_7 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_17.dl_8 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_17.u_inv_9  (.A(\u_delay_line.u_bulk_17.dl_8 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_17.dl_9 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_18.u_inv_0  (.A(\u_delay_line.bulk_17 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_18.dl_0 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_18.u_inv_1  (.A(\u_delay_line.u_bulk_18.dl_0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_18.dl_1 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_18.u_inv_10  (.A(\u_delay_line.u_bulk_18.dl_9 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_18.dl_10 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_18.u_inv_11  (.A(\u_delay_line.u_bulk_18.dl_10 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_18.dl_11 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_18.u_inv_12  (.A(\u_delay_line.u_bulk_18.dl_11 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_18.dl_12 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_18.u_inv_13  (.A(\u_delay_line.u_bulk_18.dl_12 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_18.dl_13 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_18.u_inv_14  (.A(\u_delay_line.u_bulk_18.dl_13 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_18.dl_14 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_18.u_inv_15  (.A(\u_delay_line.u_bulk_18.dl_14 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.bulk_18 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_18.u_inv_2  (.A(\u_delay_line.u_bulk_18.dl_1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_18.dl_2 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_18.u_inv_3  (.A(\u_delay_line.u_bulk_18.dl_2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_18.dl_3 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_18.u_inv_4  (.A(\u_delay_line.u_bulk_18.dl_3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_18.dl_4 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_18.u_inv_5  (.A(\u_delay_line.u_bulk_18.dl_4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_18.dl_5 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_18.u_inv_6  (.A(\u_delay_line.u_bulk_18.dl_5 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_18.dl_6 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_18.u_inv_7  (.A(\u_delay_line.u_bulk_18.dl_6 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_18.dl_7 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_18.u_inv_8  (.A(\u_delay_line.u_bulk_18.dl_7 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_18.dl_8 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_18.u_inv_9  (.A(\u_delay_line.u_bulk_18.dl_8 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_18.dl_9 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_19.u_inv_0  (.A(\u_delay_line.bulk_18 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_19.dl_0 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_19.u_inv_1  (.A(\u_delay_line.u_bulk_19.dl_0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_19.dl_1 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_19.u_inv_10  (.A(\u_delay_line.u_bulk_19.dl_9 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_19.dl_10 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_19.u_inv_11  (.A(\u_delay_line.u_bulk_19.dl_10 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_19.dl_11 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_19.u_inv_12  (.A(\u_delay_line.u_bulk_19.dl_11 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_19.dl_12 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_19.u_inv_13  (.A(\u_delay_line.u_bulk_19.dl_12 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_19.dl_13 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_19.u_inv_14  (.A(\u_delay_line.u_bulk_19.dl_13 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_19.dl_14 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_19.u_inv_15  (.A(\u_delay_line.u_bulk_19.dl_14 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.bulk_19 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_19.u_inv_2  (.A(\u_delay_line.u_bulk_19.dl_1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_19.dl_2 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_19.u_inv_3  (.A(\u_delay_line.u_bulk_19.dl_2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_19.dl_3 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_19.u_inv_4  (.A(\u_delay_line.u_bulk_19.dl_3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_19.dl_4 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_19.u_inv_5  (.A(\u_delay_line.u_bulk_19.dl_4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_19.dl_5 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_19.u_inv_6  (.A(\u_delay_line.u_bulk_19.dl_5 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_19.dl_6 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_19.u_inv_7  (.A(\u_delay_line.u_bulk_19.dl_6 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_19.dl_7 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_19.u_inv_8  (.A(\u_delay_line.u_bulk_19.dl_7 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_19.dl_8 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_19.u_inv_9  (.A(\u_delay_line.u_bulk_19.dl_8 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_19.dl_9 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_2.u_inv_0  (.A(\u_delay_line.bulk_1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_2.dl_0 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_2.u_inv_1  (.A(\u_delay_line.u_bulk_2.dl_0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_2.dl_1 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_2.u_inv_10  (.A(\u_delay_line.u_bulk_2.dl_9 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_2.dl_10 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_2.u_inv_11  (.A(\u_delay_line.u_bulk_2.dl_10 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_2.dl_11 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_2.u_inv_12  (.A(\u_delay_line.u_bulk_2.dl_11 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_2.dl_12 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_2.u_inv_13  (.A(\u_delay_line.u_bulk_2.dl_12 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_2.dl_13 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_2.u_inv_14  (.A(\u_delay_line.u_bulk_2.dl_13 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_2.dl_14 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_2.u_inv_15  (.A(\u_delay_line.u_bulk_2.dl_14 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.bulk_2 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_2.u_inv_2  (.A(\u_delay_line.u_bulk_2.dl_1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_2.dl_2 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_2.u_inv_3  (.A(\u_delay_line.u_bulk_2.dl_2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_2.dl_3 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_2.u_inv_4  (.A(\u_delay_line.u_bulk_2.dl_3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_2.dl_4 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_2.u_inv_5  (.A(\u_delay_line.u_bulk_2.dl_4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_2.dl_5 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_2.u_inv_6  (.A(\u_delay_line.u_bulk_2.dl_5 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_2.dl_6 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_2.u_inv_7  (.A(\u_delay_line.u_bulk_2.dl_6 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_2.dl_7 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_2.u_inv_8  (.A(\u_delay_line.u_bulk_2.dl_7 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_2.dl_8 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_2.u_inv_9  (.A(\u_delay_line.u_bulk_2.dl_8 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_2.dl_9 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_20.u_inv_0  (.A(\u_delay_line.bulk_19 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_20.dl_0 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_20.u_inv_1  (.A(\u_delay_line.u_bulk_20.dl_0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_20.dl_1 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_20.u_inv_10  (.A(\u_delay_line.u_bulk_20.dl_9 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_20.dl_10 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_20.u_inv_11  (.A(\u_delay_line.u_bulk_20.dl_10 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_20.dl_11 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_20.u_inv_12  (.A(\u_delay_line.u_bulk_20.dl_11 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_20.dl_12 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_20.u_inv_13  (.A(\u_delay_line.u_bulk_20.dl_12 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_20.dl_13 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_20.u_inv_14  (.A(\u_delay_line.u_bulk_20.dl_13 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_20.dl_14 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_20.u_inv_15  (.A(\u_delay_line.u_bulk_20.dl_14 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.bulk_20 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_20.u_inv_2  (.A(\u_delay_line.u_bulk_20.dl_1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_20.dl_2 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_20.u_inv_3  (.A(\u_delay_line.u_bulk_20.dl_2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_20.dl_3 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_20.u_inv_4  (.A(\u_delay_line.u_bulk_20.dl_3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_20.dl_4 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_20.u_inv_5  (.A(\u_delay_line.u_bulk_20.dl_4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_20.dl_5 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_20.u_inv_6  (.A(\u_delay_line.u_bulk_20.dl_5 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_20.dl_6 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_20.u_inv_7  (.A(\u_delay_line.u_bulk_20.dl_6 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_20.dl_7 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_20.u_inv_8  (.A(\u_delay_line.u_bulk_20.dl_7 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_20.dl_8 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_20.u_inv_9  (.A(\u_delay_line.u_bulk_20.dl_8 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_20.dl_9 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_21.u_inv_0  (.A(\u_delay_line.bulk_20 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_21.dl_0 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_21.u_inv_1  (.A(\u_delay_line.u_bulk_21.dl_0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_21.dl_1 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_21.u_inv_10  (.A(\u_delay_line.u_bulk_21.dl_9 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_21.dl_10 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_21.u_inv_11  (.A(\u_delay_line.u_bulk_21.dl_10 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_21.dl_11 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_21.u_inv_12  (.A(\u_delay_line.u_bulk_21.dl_11 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_21.dl_12 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_21.u_inv_13  (.A(\u_delay_line.u_bulk_21.dl_12 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_21.dl_13 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_21.u_inv_14  (.A(\u_delay_line.u_bulk_21.dl_13 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_21.dl_14 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_21.u_inv_15  (.A(\u_delay_line.u_bulk_21.dl_14 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.dl_0 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_21.u_inv_2  (.A(\u_delay_line.u_bulk_21.dl_1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_21.dl_2 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_21.u_inv_3  (.A(\u_delay_line.u_bulk_21.dl_2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_21.dl_3 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_21.u_inv_4  (.A(\u_delay_line.u_bulk_21.dl_3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_21.dl_4 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_21.u_inv_5  (.A(\u_delay_line.u_bulk_21.dl_4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_21.dl_5 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_21.u_inv_6  (.A(\u_delay_line.u_bulk_21.dl_5 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_21.dl_6 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_21.u_inv_7  (.A(\u_delay_line.u_bulk_21.dl_6 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_21.dl_7 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_21.u_inv_8  (.A(\u_delay_line.u_bulk_21.dl_7 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_21.dl_8 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_21.u_inv_9  (.A(\u_delay_line.u_bulk_21.dl_8 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_21.dl_9 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_3.u_inv_0  (.A(\u_delay_line.bulk_2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_3.dl_0 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_3.u_inv_1  (.A(\u_delay_line.u_bulk_3.dl_0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_3.dl_1 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_3.u_inv_10  (.A(\u_delay_line.u_bulk_3.dl_9 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_3.dl_10 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_3.u_inv_11  (.A(\u_delay_line.u_bulk_3.dl_10 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_3.dl_11 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_3.u_inv_12  (.A(\u_delay_line.u_bulk_3.dl_11 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_3.dl_12 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_3.u_inv_13  (.A(\u_delay_line.u_bulk_3.dl_12 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_3.dl_13 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_3.u_inv_14  (.A(\u_delay_line.u_bulk_3.dl_13 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_3.dl_14 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_3.u_inv_15  (.A(\u_delay_line.u_bulk_3.dl_14 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.bulk_3 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_3.u_inv_2  (.A(\u_delay_line.u_bulk_3.dl_1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_3.dl_2 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_3.u_inv_3  (.A(\u_delay_line.u_bulk_3.dl_2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_3.dl_3 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_3.u_inv_4  (.A(\u_delay_line.u_bulk_3.dl_3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_3.dl_4 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_3.u_inv_5  (.A(\u_delay_line.u_bulk_3.dl_4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_3.dl_5 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_3.u_inv_6  (.A(\u_delay_line.u_bulk_3.dl_5 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_3.dl_6 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_3.u_inv_7  (.A(\u_delay_line.u_bulk_3.dl_6 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_3.dl_7 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_3.u_inv_8  (.A(\u_delay_line.u_bulk_3.dl_7 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_3.dl_8 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_3.u_inv_9  (.A(\u_delay_line.u_bulk_3.dl_8 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_3.dl_9 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_4.u_inv_0  (.A(\u_delay_line.bulk_3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_4.dl_0 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_4.u_inv_1  (.A(\u_delay_line.u_bulk_4.dl_0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_4.dl_1 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_4.u_inv_10  (.A(\u_delay_line.u_bulk_4.dl_9 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_4.dl_10 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_4.u_inv_11  (.A(\u_delay_line.u_bulk_4.dl_10 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_4.dl_11 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_4.u_inv_12  (.A(\u_delay_line.u_bulk_4.dl_11 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_4.dl_12 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_4.u_inv_13  (.A(\u_delay_line.u_bulk_4.dl_12 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_4.dl_13 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_4.u_inv_14  (.A(\u_delay_line.u_bulk_4.dl_13 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_4.dl_14 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_4.u_inv_15  (.A(\u_delay_line.u_bulk_4.dl_14 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.bulk_4 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_4.u_inv_2  (.A(\u_delay_line.u_bulk_4.dl_1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_4.dl_2 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_4.u_inv_3  (.A(\u_delay_line.u_bulk_4.dl_2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_4.dl_3 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_4.u_inv_4  (.A(\u_delay_line.u_bulk_4.dl_3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_4.dl_4 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_4.u_inv_5  (.A(\u_delay_line.u_bulk_4.dl_4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_4.dl_5 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_4.u_inv_6  (.A(\u_delay_line.u_bulk_4.dl_5 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_4.dl_6 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_4.u_inv_7  (.A(\u_delay_line.u_bulk_4.dl_6 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_4.dl_7 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_4.u_inv_8  (.A(\u_delay_line.u_bulk_4.dl_7 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_4.dl_8 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_4.u_inv_9  (.A(\u_delay_line.u_bulk_4.dl_8 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_4.dl_9 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_5.u_inv_0  (.A(\u_delay_line.bulk_4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_5.dl_0 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_5.u_inv_1  (.A(\u_delay_line.u_bulk_5.dl_0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_5.dl_1 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_5.u_inv_10  (.A(\u_delay_line.u_bulk_5.dl_9 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_5.dl_10 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_5.u_inv_11  (.A(\u_delay_line.u_bulk_5.dl_10 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_5.dl_11 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_5.u_inv_12  (.A(\u_delay_line.u_bulk_5.dl_11 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_5.dl_12 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_5.u_inv_13  (.A(\u_delay_line.u_bulk_5.dl_12 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_5.dl_13 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_5.u_inv_14  (.A(\u_delay_line.u_bulk_5.dl_13 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_5.dl_14 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_5.u_inv_15  (.A(\u_delay_line.u_bulk_5.dl_14 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.bulk_5 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_5.u_inv_2  (.A(\u_delay_line.u_bulk_5.dl_1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_5.dl_2 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_5.u_inv_3  (.A(\u_delay_line.u_bulk_5.dl_2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_5.dl_3 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_5.u_inv_4  (.A(\u_delay_line.u_bulk_5.dl_3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_5.dl_4 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_5.u_inv_5  (.A(\u_delay_line.u_bulk_5.dl_4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_5.dl_5 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_5.u_inv_6  (.A(\u_delay_line.u_bulk_5.dl_5 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_5.dl_6 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_5.u_inv_7  (.A(\u_delay_line.u_bulk_5.dl_6 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_5.dl_7 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_5.u_inv_8  (.A(\u_delay_line.u_bulk_5.dl_7 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_5.dl_8 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_5.u_inv_9  (.A(\u_delay_line.u_bulk_5.dl_8 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_5.dl_9 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_6.u_inv_0  (.A(\u_delay_line.bulk_5 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_6.dl_0 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_6.u_inv_1  (.A(\u_delay_line.u_bulk_6.dl_0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_6.dl_1 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_6.u_inv_10  (.A(\u_delay_line.u_bulk_6.dl_9 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_6.dl_10 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_6.u_inv_11  (.A(\u_delay_line.u_bulk_6.dl_10 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_6.dl_11 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_6.u_inv_12  (.A(\u_delay_line.u_bulk_6.dl_11 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_6.dl_12 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_6.u_inv_13  (.A(\u_delay_line.u_bulk_6.dl_12 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_6.dl_13 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_6.u_inv_14  (.A(\u_delay_line.u_bulk_6.dl_13 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_6.dl_14 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_6.u_inv_15  (.A(\u_delay_line.u_bulk_6.dl_14 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.bulk_6 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_6.u_inv_2  (.A(\u_delay_line.u_bulk_6.dl_1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_6.dl_2 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_6.u_inv_3  (.A(\u_delay_line.u_bulk_6.dl_2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_6.dl_3 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_6.u_inv_4  (.A(\u_delay_line.u_bulk_6.dl_3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_6.dl_4 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_6.u_inv_5  (.A(\u_delay_line.u_bulk_6.dl_4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_6.dl_5 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_6.u_inv_6  (.A(\u_delay_line.u_bulk_6.dl_5 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_6.dl_6 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_6.u_inv_7  (.A(\u_delay_line.u_bulk_6.dl_6 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_6.dl_7 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_6.u_inv_8  (.A(\u_delay_line.u_bulk_6.dl_7 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_6.dl_8 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_6.u_inv_9  (.A(\u_delay_line.u_bulk_6.dl_8 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_6.dl_9 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_7.u_inv_0  (.A(\u_delay_line.bulk_6 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_7.dl_0 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_7.u_inv_1  (.A(\u_delay_line.u_bulk_7.dl_0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_7.dl_1 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_7.u_inv_10  (.A(\u_delay_line.u_bulk_7.dl_9 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_7.dl_10 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_7.u_inv_11  (.A(\u_delay_line.u_bulk_7.dl_10 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_7.dl_11 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_7.u_inv_12  (.A(\u_delay_line.u_bulk_7.dl_11 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_7.dl_12 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_7.u_inv_13  (.A(\u_delay_line.u_bulk_7.dl_12 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_7.dl_13 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_7.u_inv_14  (.A(\u_delay_line.u_bulk_7.dl_13 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_7.dl_14 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_7.u_inv_15  (.A(\u_delay_line.u_bulk_7.dl_14 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.bulk_7 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_7.u_inv_2  (.A(\u_delay_line.u_bulk_7.dl_1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_7.dl_2 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_7.u_inv_3  (.A(\u_delay_line.u_bulk_7.dl_2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_7.dl_3 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_7.u_inv_4  (.A(\u_delay_line.u_bulk_7.dl_3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_7.dl_4 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_7.u_inv_5  (.A(\u_delay_line.u_bulk_7.dl_4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_7.dl_5 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_7.u_inv_6  (.A(\u_delay_line.u_bulk_7.dl_5 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_7.dl_6 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_7.u_inv_7  (.A(\u_delay_line.u_bulk_7.dl_6 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_7.dl_7 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_7.u_inv_8  (.A(\u_delay_line.u_bulk_7.dl_7 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_7.dl_8 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_7.u_inv_9  (.A(\u_delay_line.u_bulk_7.dl_8 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_7.dl_9 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_8.u_inv_0  (.A(\u_delay_line.bulk_7 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_8.dl_0 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_8.u_inv_1  (.A(\u_delay_line.u_bulk_8.dl_0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_8.dl_1 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_8.u_inv_10  (.A(\u_delay_line.u_bulk_8.dl_9 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_8.dl_10 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_8.u_inv_11  (.A(\u_delay_line.u_bulk_8.dl_10 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_8.dl_11 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_8.u_inv_12  (.A(\u_delay_line.u_bulk_8.dl_11 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_8.dl_12 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_8.u_inv_13  (.A(\u_delay_line.u_bulk_8.dl_12 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_8.dl_13 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_8.u_inv_14  (.A(\u_delay_line.u_bulk_8.dl_13 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_8.dl_14 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_8.u_inv_15  (.A(\u_delay_line.u_bulk_8.dl_14 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.bulk_8 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_8.u_inv_2  (.A(\u_delay_line.u_bulk_8.dl_1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_8.dl_2 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_8.u_inv_3  (.A(\u_delay_line.u_bulk_8.dl_2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_8.dl_3 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_8.u_inv_4  (.A(\u_delay_line.u_bulk_8.dl_3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_8.dl_4 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_8.u_inv_5  (.A(\u_delay_line.u_bulk_8.dl_4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_8.dl_5 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_8.u_inv_6  (.A(\u_delay_line.u_bulk_8.dl_5 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_8.dl_6 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_8.u_inv_7  (.A(\u_delay_line.u_bulk_8.dl_6 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_8.dl_7 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_8.u_inv_8  (.A(\u_delay_line.u_bulk_8.dl_7 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_8.dl_8 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_8.u_inv_9  (.A(\u_delay_line.u_bulk_8.dl_8 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_8.dl_9 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_9.u_inv_0  (.A(\u_delay_line.bulk_8 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_9.dl_0 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_9.u_inv_1  (.A(\u_delay_line.u_bulk_9.dl_0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_9.dl_1 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_9.u_inv_10  (.A(\u_delay_line.u_bulk_9.dl_9 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_9.dl_10 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_9.u_inv_11  (.A(\u_delay_line.u_bulk_9.dl_10 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_9.dl_11 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_9.u_inv_12  (.A(\u_delay_line.u_bulk_9.dl_11 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_9.dl_12 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_9.u_inv_13  (.A(\u_delay_line.u_bulk_9.dl_12 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_9.dl_13 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_9.u_inv_14  (.A(\u_delay_line.u_bulk_9.dl_13 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_9.dl_14 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_9.u_inv_15  (.A(\u_delay_line.u_bulk_9.dl_14 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.bulk_9 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_9.u_inv_2  (.A(\u_delay_line.u_bulk_9.dl_1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_9.dl_2 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_9.u_inv_3  (.A(\u_delay_line.u_bulk_9.dl_2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_9.dl_3 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_9.u_inv_4  (.A(\u_delay_line.u_bulk_9.dl_3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_9.dl_4 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_9.u_inv_5  (.A(\u_delay_line.u_bulk_9.dl_4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_9.dl_5 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_9.u_inv_6  (.A(\u_delay_line.u_bulk_9.dl_5 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_9.dl_6 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_9.u_inv_7  (.A(\u_delay_line.u_bulk_9.dl_6 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_9.dl_7 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_9.u_inv_8  (.A(\u_delay_line.u_bulk_9.dl_7 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_9.dl_8 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_bulk_9.u_inv_9  (.A(\u_delay_line.u_bulk_9.dl_8 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_bulk_9.dl_9 ));
 sky130_fd_sc_hd__dfrtp_1 \u_delay_line.u_dl_0.u_ff  (.CLK(clknet_4_1_0_clk),
    .D(\u_delay_line.dl_1 ),
    .RESET_B(net4),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\u_delay_line.data_0 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_0.u_inv_0  (.A(\u_delay_line.dl_0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_0.dl_0 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_0.u_inv_1  (.A(\u_delay_line.u_dl_0.dl_0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_0.dl_1 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_0.u_inv_10  (.A(\u_delay_line.u_dl_0.dl_9 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_0.dl_10 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_0.u_inv_11  (.A(\u_delay_line.u_dl_0.dl_10 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.dl_1 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_0.u_inv_2  (.A(\u_delay_line.u_dl_0.dl_1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_0.dl_2 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_0.u_inv_3  (.A(\u_delay_line.u_dl_0.dl_2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_0.dl_3 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_0.u_inv_4  (.A(\u_delay_line.u_dl_0.dl_3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_0.dl_4 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_0.u_inv_5  (.A(\u_delay_line.u_dl_0.dl_4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_0.dl_5 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_0.u_inv_6  (.A(\u_delay_line.u_dl_0.dl_5 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_0.dl_6 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_0.u_inv_7  (.A(\u_delay_line.u_dl_0.dl_6 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_0.dl_7 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_0.u_inv_8  (.A(\u_delay_line.u_dl_0.dl_7 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_0.dl_8 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_0.u_inv_9  (.A(\u_delay_line.u_dl_0.dl_8 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_0.dl_9 ));
 sky130_fd_sc_hd__dfrtp_1 \u_delay_line.u_dl_1.u_ff  (.CLK(clknet_4_1_0_clk),
    .D(\u_delay_line.dl_2 ),
    .RESET_B(net4),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\u_delay_line.data_1 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_1.u_inv_0  (.A(\u_delay_line.dl_1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_1.dl_0 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_1.u_inv_1  (.A(\u_delay_line.u_dl_1.dl_0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_1.dl_1 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_1.u_inv_10  (.A(\u_delay_line.u_dl_1.dl_9 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_1.dl_10 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_1.u_inv_11  (.A(\u_delay_line.u_dl_1.dl_10 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.dl_2 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_1.u_inv_2  (.A(\u_delay_line.u_dl_1.dl_1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_1.dl_2 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_1.u_inv_3  (.A(\u_delay_line.u_dl_1.dl_2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_1.dl_3 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_1.u_inv_4  (.A(\u_delay_line.u_dl_1.dl_3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_1.dl_4 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_1.u_inv_5  (.A(\u_delay_line.u_dl_1.dl_4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_1.dl_5 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_1.u_inv_6  (.A(\u_delay_line.u_dl_1.dl_5 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_1.dl_6 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_1.u_inv_7  (.A(\u_delay_line.u_dl_1.dl_6 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_1.dl_7 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_1.u_inv_8  (.A(\u_delay_line.u_dl_1.dl_7 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_1.dl_8 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_1.u_inv_9  (.A(\u_delay_line.u_dl_1.dl_8 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_1.dl_9 ));
 sky130_fd_sc_hd__dfrtp_1 \u_delay_line.u_dl_10.u_ff  (.CLK(clknet_4_4_0_clk),
    .D(\u_delay_line.dl_11 ),
    .RESET_B(net7),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\u_delay_line.data_10 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_10.u_inv_0  (.A(\u_delay_line.dl_10 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_10.dl_0 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_10.u_inv_1  (.A(\u_delay_line.u_dl_10.dl_0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_10.dl_1 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_10.u_inv_10  (.A(\u_delay_line.u_dl_10.dl_9 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_10.dl_10 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_10.u_inv_11  (.A(\u_delay_line.u_dl_10.dl_10 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.dl_11 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_10.u_inv_2  (.A(\u_delay_line.u_dl_10.dl_1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_10.dl_2 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_10.u_inv_3  (.A(\u_delay_line.u_dl_10.dl_2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_10.dl_3 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_10.u_inv_4  (.A(\u_delay_line.u_dl_10.dl_3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_10.dl_4 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_10.u_inv_5  (.A(\u_delay_line.u_dl_10.dl_4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_10.dl_5 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_10.u_inv_6  (.A(\u_delay_line.u_dl_10.dl_5 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_10.dl_6 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_10.u_inv_7  (.A(\u_delay_line.u_dl_10.dl_6 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_10.dl_7 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_10.u_inv_8  (.A(\u_delay_line.u_dl_10.dl_7 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_10.dl_8 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_10.u_inv_9  (.A(\u_delay_line.u_dl_10.dl_8 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_10.dl_9 ));
 sky130_fd_sc_hd__dfrtp_1 \u_delay_line.u_dl_11.u_ff  (.CLK(clknet_4_5_0_clk),
    .D(\u_delay_line.dl_12 ),
    .RESET_B(net7),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\u_delay_line.data_11 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_11.u_inv_0  (.A(\u_delay_line.dl_11 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_11.dl_0 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_11.u_inv_1  (.A(\u_delay_line.u_dl_11.dl_0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_11.dl_1 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_11.u_inv_10  (.A(\u_delay_line.u_dl_11.dl_9 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_11.dl_10 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_11.u_inv_11  (.A(\u_delay_line.u_dl_11.dl_10 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.dl_12 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_11.u_inv_2  (.A(\u_delay_line.u_dl_11.dl_1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_11.dl_2 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_11.u_inv_3  (.A(\u_delay_line.u_dl_11.dl_2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_11.dl_3 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_11.u_inv_4  (.A(\u_delay_line.u_dl_11.dl_3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_11.dl_4 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_11.u_inv_5  (.A(\u_delay_line.u_dl_11.dl_4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_11.dl_5 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_11.u_inv_6  (.A(\u_delay_line.u_dl_11.dl_5 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_11.dl_6 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_11.u_inv_7  (.A(\u_delay_line.u_dl_11.dl_6 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_11.dl_7 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_11.u_inv_8  (.A(\u_delay_line.u_dl_11.dl_7 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_11.dl_8 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_11.u_inv_9  (.A(\u_delay_line.u_dl_11.dl_8 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_11.dl_9 ));
 sky130_fd_sc_hd__dfrtp_1 \u_delay_line.u_dl_12.u_ff  (.CLK(clknet_4_5_0_clk),
    .D(\u_delay_line.dl_13 ),
    .RESET_B(net10),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\u_delay_line.data_12 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_12.u_inv_0  (.A(\u_delay_line.dl_12 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_12.dl_0 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_12.u_inv_1  (.A(\u_delay_line.u_dl_12.dl_0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_12.dl_1 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_12.u_inv_10  (.A(\u_delay_line.u_dl_12.dl_9 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_12.dl_10 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_12.u_inv_11  (.A(\u_delay_line.u_dl_12.dl_10 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.dl_13 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_12.u_inv_2  (.A(\u_delay_line.u_dl_12.dl_1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_12.dl_2 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_12.u_inv_3  (.A(\u_delay_line.u_dl_12.dl_2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_12.dl_3 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_12.u_inv_4  (.A(\u_delay_line.u_dl_12.dl_3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_12.dl_4 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_12.u_inv_5  (.A(\u_delay_line.u_dl_12.dl_4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_12.dl_5 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_12.u_inv_6  (.A(\u_delay_line.u_dl_12.dl_5 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_12.dl_6 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_12.u_inv_7  (.A(\u_delay_line.u_dl_12.dl_6 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_12.dl_7 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_12.u_inv_8  (.A(\u_delay_line.u_dl_12.dl_7 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_12.dl_8 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_12.u_inv_9  (.A(\u_delay_line.u_dl_12.dl_8 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_12.dl_9 ));
 sky130_fd_sc_hd__dfrtp_1 \u_delay_line.u_dl_13.u_ff  (.CLK(clknet_4_5_0_clk),
    .D(\u_delay_line.dl_14 ),
    .RESET_B(net9),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\u_delay_line.data_13 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_13.u_inv_0  (.A(\u_delay_line.dl_13 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_13.dl_0 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_13.u_inv_1  (.A(\u_delay_line.u_dl_13.dl_0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_13.dl_1 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_13.u_inv_10  (.A(\u_delay_line.u_dl_13.dl_9 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_13.dl_10 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_13.u_inv_11  (.A(\u_delay_line.u_dl_13.dl_10 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.dl_14 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_13.u_inv_2  (.A(\u_delay_line.u_dl_13.dl_1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_13.dl_2 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_13.u_inv_3  (.A(\u_delay_line.u_dl_13.dl_2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_13.dl_3 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_13.u_inv_4  (.A(\u_delay_line.u_dl_13.dl_3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_13.dl_4 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_13.u_inv_5  (.A(\u_delay_line.u_dl_13.dl_4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_13.dl_5 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_13.u_inv_6  (.A(\u_delay_line.u_dl_13.dl_5 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_13.dl_6 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_13.u_inv_7  (.A(\u_delay_line.u_dl_13.dl_6 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_13.dl_7 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_13.u_inv_8  (.A(\u_delay_line.u_dl_13.dl_7 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_13.dl_8 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_13.u_inv_9  (.A(\u_delay_line.u_dl_13.dl_8 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_13.dl_9 ));
 sky130_fd_sc_hd__dfrtp_1 \u_delay_line.u_dl_14.u_ff  (.CLK(clknet_4_4_0_clk),
    .D(\u_delay_line.dl_15 ),
    .RESET_B(net7),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\u_delay_line.data_14 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_14.u_inv_0  (.A(\u_delay_line.dl_14 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_14.dl_0 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_14.u_inv_1  (.A(\u_delay_line.u_dl_14.dl_0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_14.dl_1 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_14.u_inv_10  (.A(\u_delay_line.u_dl_14.dl_9 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_14.dl_10 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_14.u_inv_11  (.A(\u_delay_line.u_dl_14.dl_10 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.dl_15 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_14.u_inv_2  (.A(\u_delay_line.u_dl_14.dl_1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_14.dl_2 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_14.u_inv_3  (.A(\u_delay_line.u_dl_14.dl_2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_14.dl_3 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_14.u_inv_4  (.A(\u_delay_line.u_dl_14.dl_3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_14.dl_4 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_14.u_inv_5  (.A(\u_delay_line.u_dl_14.dl_4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_14.dl_5 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_14.u_inv_6  (.A(\u_delay_line.u_dl_14.dl_5 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_14.dl_6 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_14.u_inv_7  (.A(\u_delay_line.u_dl_14.dl_6 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_14.dl_7 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_14.u_inv_8  (.A(\u_delay_line.u_dl_14.dl_7 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_14.dl_8 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_14.u_inv_9  (.A(\u_delay_line.u_dl_14.dl_8 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_14.dl_9 ));
 sky130_fd_sc_hd__dfrtp_1 \u_delay_line.u_dl_15.u_ff  (.CLK(clknet_4_6_0_clk),
    .D(\u_delay_line.dl_16 ),
    .RESET_B(net8),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\u_delay_line.data_15 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_15.u_inv_0  (.A(\u_delay_line.dl_15 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_15.dl_0 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_15.u_inv_1  (.A(\u_delay_line.u_dl_15.dl_0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_15.dl_1 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_15.u_inv_10  (.A(\u_delay_line.u_dl_15.dl_9 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_15.dl_10 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_15.u_inv_11  (.A(\u_delay_line.u_dl_15.dl_10 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.dl_16 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_15.u_inv_2  (.A(\u_delay_line.u_dl_15.dl_1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_15.dl_2 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_15.u_inv_3  (.A(\u_delay_line.u_dl_15.dl_2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_15.dl_3 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_15.u_inv_4  (.A(\u_delay_line.u_dl_15.dl_3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_15.dl_4 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_15.u_inv_5  (.A(\u_delay_line.u_dl_15.dl_4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_15.dl_5 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_15.u_inv_6  (.A(\u_delay_line.u_dl_15.dl_5 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_15.dl_6 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_15.u_inv_7  (.A(\u_delay_line.u_dl_15.dl_6 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_15.dl_7 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_15.u_inv_8  (.A(\u_delay_line.u_dl_15.dl_7 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_15.dl_8 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_15.u_inv_9  (.A(\u_delay_line.u_dl_15.dl_8 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_15.dl_9 ));
 sky130_fd_sc_hd__dfrtp_1 \u_delay_line.u_dl_16.u_ff  (.CLK(clknet_4_4_0_clk),
    .D(\u_delay_line.dl_17 ),
    .RESET_B(net7),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\u_delay_line.data_16 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_16.u_inv_0  (.A(\u_delay_line.dl_16 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_16.dl_0 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_16.u_inv_1  (.A(\u_delay_line.u_dl_16.dl_0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_16.dl_1 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_16.u_inv_10  (.A(\u_delay_line.u_dl_16.dl_9 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_16.dl_10 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_16.u_inv_11  (.A(\u_delay_line.u_dl_16.dl_10 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.dl_17 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_16.u_inv_2  (.A(\u_delay_line.u_dl_16.dl_1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_16.dl_2 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_16.u_inv_3  (.A(\u_delay_line.u_dl_16.dl_2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_16.dl_3 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_16.u_inv_4  (.A(\u_delay_line.u_dl_16.dl_3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_16.dl_4 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_16.u_inv_5  (.A(\u_delay_line.u_dl_16.dl_4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_16.dl_5 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_16.u_inv_6  (.A(\u_delay_line.u_dl_16.dl_5 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_16.dl_6 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_16.u_inv_7  (.A(\u_delay_line.u_dl_16.dl_6 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_16.dl_7 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_16.u_inv_8  (.A(\u_delay_line.u_dl_16.dl_7 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_16.dl_8 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_16.u_inv_9  (.A(\u_delay_line.u_dl_16.dl_8 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_16.dl_9 ));
 sky130_fd_sc_hd__dfrtp_1 \u_delay_line.u_dl_17.u_ff  (.CLK(clknet_4_4_0_clk),
    .D(\u_delay_line.dl_18 ),
    .RESET_B(net7),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\u_delay_line.data_17 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_17.u_inv_0  (.A(\u_delay_line.dl_17 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_17.dl_0 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_17.u_inv_1  (.A(\u_delay_line.u_dl_17.dl_0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_17.dl_1 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_17.u_inv_10  (.A(\u_delay_line.u_dl_17.dl_9 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_17.dl_10 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_17.u_inv_11  (.A(\u_delay_line.u_dl_17.dl_10 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.dl_18 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_17.u_inv_2  (.A(\u_delay_line.u_dl_17.dl_1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_17.dl_2 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_17.u_inv_3  (.A(\u_delay_line.u_dl_17.dl_2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_17.dl_3 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_17.u_inv_4  (.A(\u_delay_line.u_dl_17.dl_3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_17.dl_4 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_17.u_inv_5  (.A(\u_delay_line.u_dl_17.dl_4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_17.dl_5 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_17.u_inv_6  (.A(\u_delay_line.u_dl_17.dl_5 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_17.dl_6 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_17.u_inv_7  (.A(\u_delay_line.u_dl_17.dl_6 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_17.dl_7 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_17.u_inv_8  (.A(\u_delay_line.u_dl_17.dl_7 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_17.dl_8 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_17.u_inv_9  (.A(\u_delay_line.u_dl_17.dl_8 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_17.dl_9 ));
 sky130_fd_sc_hd__dfrtp_1 \u_delay_line.u_dl_18.u_ff  (.CLK(clknet_4_1_0_clk),
    .D(\u_delay_line.dl_19 ),
    .RESET_B(net4),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\u_delay_line.data_18 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_18.u_inv_0  (.A(\u_delay_line.dl_18 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_18.dl_0 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_18.u_inv_1  (.A(\u_delay_line.u_dl_18.dl_0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_18.dl_1 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_18.u_inv_10  (.A(\u_delay_line.u_dl_18.dl_9 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_18.dl_10 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_18.u_inv_11  (.A(\u_delay_line.u_dl_18.dl_10 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.dl_19 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_18.u_inv_2  (.A(\u_delay_line.u_dl_18.dl_1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_18.dl_2 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_18.u_inv_3  (.A(\u_delay_line.u_dl_18.dl_2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_18.dl_3 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_18.u_inv_4  (.A(\u_delay_line.u_dl_18.dl_3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_18.dl_4 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_18.u_inv_5  (.A(\u_delay_line.u_dl_18.dl_4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_18.dl_5 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_18.u_inv_6  (.A(\u_delay_line.u_dl_18.dl_5 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_18.dl_6 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_18.u_inv_7  (.A(\u_delay_line.u_dl_18.dl_6 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_18.dl_7 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_18.u_inv_8  (.A(\u_delay_line.u_dl_18.dl_7 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_18.dl_8 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_18.u_inv_9  (.A(\u_delay_line.u_dl_18.dl_8 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_18.dl_9 ));
 sky130_fd_sc_hd__dfrtp_1 \u_delay_line.u_dl_19.u_ff  (.CLK(clknet_4_0_0_clk),
    .D(\u_delay_line.dl_20 ),
    .RESET_B(net3),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\u_delay_line.data_19 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_19.u_inv_0  (.A(\u_delay_line.dl_19 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_19.dl_0 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_19.u_inv_1  (.A(\u_delay_line.u_dl_19.dl_0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_19.dl_1 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_19.u_inv_10  (.A(\u_delay_line.u_dl_19.dl_9 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_19.dl_10 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_19.u_inv_11  (.A(\u_delay_line.u_dl_19.dl_10 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.dl_20 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_19.u_inv_2  (.A(\u_delay_line.u_dl_19.dl_1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_19.dl_2 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_19.u_inv_3  (.A(\u_delay_line.u_dl_19.dl_2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_19.dl_3 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_19.u_inv_4  (.A(\u_delay_line.u_dl_19.dl_3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_19.dl_4 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_19.u_inv_5  (.A(\u_delay_line.u_dl_19.dl_4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_19.dl_5 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_19.u_inv_6  (.A(\u_delay_line.u_dl_19.dl_5 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_19.dl_6 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_19.u_inv_7  (.A(\u_delay_line.u_dl_19.dl_6 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_19.dl_7 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_19.u_inv_8  (.A(\u_delay_line.u_dl_19.dl_7 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_19.dl_8 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_19.u_inv_9  (.A(\u_delay_line.u_dl_19.dl_8 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_19.dl_9 ));
 sky130_fd_sc_hd__dfrtp_1 \u_delay_line.u_dl_2.u_ff  (.CLK(clknet_4_0_0_clk),
    .D(\u_delay_line.dl_3 ),
    .RESET_B(net3),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\u_delay_line.data_2 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_2.u_inv_0  (.A(\u_delay_line.dl_2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_2.dl_0 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_2.u_inv_1  (.A(\u_delay_line.u_dl_2.dl_0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_2.dl_1 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_2.u_inv_10  (.A(\u_delay_line.u_dl_2.dl_9 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_2.dl_10 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_2.u_inv_11  (.A(\u_delay_line.u_dl_2.dl_10 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.dl_3 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_2.u_inv_2  (.A(\u_delay_line.u_dl_2.dl_1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_2.dl_2 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_2.u_inv_3  (.A(\u_delay_line.u_dl_2.dl_2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_2.dl_3 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_2.u_inv_4  (.A(\u_delay_line.u_dl_2.dl_3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_2.dl_4 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_2.u_inv_5  (.A(\u_delay_line.u_dl_2.dl_4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_2.dl_5 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_2.u_inv_6  (.A(\u_delay_line.u_dl_2.dl_5 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_2.dl_6 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_2.u_inv_7  (.A(\u_delay_line.u_dl_2.dl_6 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_2.dl_7 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_2.u_inv_8  (.A(\u_delay_line.u_dl_2.dl_7 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_2.dl_8 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_2.u_inv_9  (.A(\u_delay_line.u_dl_2.dl_8 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_2.dl_9 ));
 sky130_fd_sc_hd__dfrtp_1 \u_delay_line.u_dl_20.u_ff  (.CLK(clknet_4_0_0_clk),
    .D(\u_delay_line.dl_21 ),
    .RESET_B(net3),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\u_delay_line.data_20 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_20.u_inv_0  (.A(\u_delay_line.dl_20 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_20.dl_0 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_20.u_inv_1  (.A(\u_delay_line.u_dl_20.dl_0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_20.dl_1 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_20.u_inv_10  (.A(\u_delay_line.u_dl_20.dl_9 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_20.dl_10 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_20.u_inv_11  (.A(\u_delay_line.u_dl_20.dl_10 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.dl_21 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_20.u_inv_2  (.A(\u_delay_line.u_dl_20.dl_1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_20.dl_2 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_20.u_inv_3  (.A(\u_delay_line.u_dl_20.dl_2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_20.dl_3 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_20.u_inv_4  (.A(\u_delay_line.u_dl_20.dl_3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_20.dl_4 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_20.u_inv_5  (.A(\u_delay_line.u_dl_20.dl_4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_20.dl_5 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_20.u_inv_6  (.A(\u_delay_line.u_dl_20.dl_5 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_20.dl_6 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_20.u_inv_7  (.A(\u_delay_line.u_dl_20.dl_6 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_20.dl_7 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_20.u_inv_8  (.A(\u_delay_line.u_dl_20.dl_7 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_20.dl_8 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_20.u_inv_9  (.A(\u_delay_line.u_dl_20.dl_8 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_20.dl_9 ));
 sky130_fd_sc_hd__dfrtp_1 \u_delay_line.u_dl_21.u_ff  (.CLK(clknet_4_0_0_clk),
    .D(\u_delay_line.dl_22 ),
    .RESET_B(net3),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\u_delay_line.data_21 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_21.u_inv_0  (.A(\u_delay_line.dl_21 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_21.dl_0 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_21.u_inv_1  (.A(\u_delay_line.u_dl_21.dl_0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_21.dl_1 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_21.u_inv_10  (.A(\u_delay_line.u_dl_21.dl_9 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_21.dl_10 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_21.u_inv_11  (.A(\u_delay_line.u_dl_21.dl_10 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.dl_22 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_21.u_inv_2  (.A(\u_delay_line.u_dl_21.dl_1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_21.dl_2 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_21.u_inv_3  (.A(\u_delay_line.u_dl_21.dl_2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_21.dl_3 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_21.u_inv_4  (.A(\u_delay_line.u_dl_21.dl_3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_21.dl_4 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_21.u_inv_5  (.A(\u_delay_line.u_dl_21.dl_4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_21.dl_5 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_21.u_inv_6  (.A(\u_delay_line.u_dl_21.dl_5 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_21.dl_6 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_21.u_inv_7  (.A(\u_delay_line.u_dl_21.dl_6 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_21.dl_7 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_21.u_inv_8  (.A(\u_delay_line.u_dl_21.dl_7 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_21.dl_8 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_21.u_inv_9  (.A(\u_delay_line.u_dl_21.dl_8 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_21.dl_9 ));
 sky130_fd_sc_hd__dfrtp_1 \u_delay_line.u_dl_22.u_ff  (.CLK(clknet_4_0_0_clk),
    .D(\u_delay_line.dl_23 ),
    .RESET_B(net3),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\u_delay_line.data_22 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_22.u_inv_0  (.A(\u_delay_line.dl_22 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_22.dl_0 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_22.u_inv_1  (.A(\u_delay_line.u_dl_22.dl_0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_22.dl_1 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_22.u_inv_10  (.A(\u_delay_line.u_dl_22.dl_9 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_22.dl_10 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_22.u_inv_11  (.A(\u_delay_line.u_dl_22.dl_10 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.dl_23 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_22.u_inv_2  (.A(\u_delay_line.u_dl_22.dl_1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_22.dl_2 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_22.u_inv_3  (.A(\u_delay_line.u_dl_22.dl_2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_22.dl_3 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_22.u_inv_4  (.A(\u_delay_line.u_dl_22.dl_3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_22.dl_4 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_22.u_inv_5  (.A(\u_delay_line.u_dl_22.dl_4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_22.dl_5 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_22.u_inv_6  (.A(\u_delay_line.u_dl_22.dl_5 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_22.dl_6 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_22.u_inv_7  (.A(\u_delay_line.u_dl_22.dl_6 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_22.dl_7 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_22.u_inv_8  (.A(\u_delay_line.u_dl_22.dl_7 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_22.dl_8 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_22.u_inv_9  (.A(\u_delay_line.u_dl_22.dl_8 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_22.dl_9 ));
 sky130_fd_sc_hd__dfrtp_1 \u_delay_line.u_dl_23.u_ff  (.CLK(clknet_4_0_0_clk),
    .D(\u_delay_line.dl_24 ),
    .RESET_B(net5),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\u_delay_line.data_23 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_23.u_inv_0  (.A(\u_delay_line.dl_23 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_23.dl_0 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_23.u_inv_1  (.A(\u_delay_line.u_dl_23.dl_0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_23.dl_1 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_23.u_inv_10  (.A(\u_delay_line.u_dl_23.dl_9 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_23.dl_10 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_23.u_inv_11  (.A(\u_delay_line.u_dl_23.dl_10 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.dl_24 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_23.u_inv_2  (.A(\u_delay_line.u_dl_23.dl_1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_23.dl_2 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_23.u_inv_3  (.A(\u_delay_line.u_dl_23.dl_2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_23.dl_3 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_23.u_inv_4  (.A(\u_delay_line.u_dl_23.dl_3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_23.dl_4 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_23.u_inv_5  (.A(\u_delay_line.u_dl_23.dl_4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_23.dl_5 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_23.u_inv_6  (.A(\u_delay_line.u_dl_23.dl_5 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_23.dl_6 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_23.u_inv_7  (.A(\u_delay_line.u_dl_23.dl_6 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_23.dl_7 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_23.u_inv_8  (.A(\u_delay_line.u_dl_23.dl_7 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_23.dl_8 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_23.u_inv_9  (.A(\u_delay_line.u_dl_23.dl_8 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_23.dl_9 ));
 sky130_fd_sc_hd__dfrtp_1 \u_delay_line.u_dl_24.u_ff  (.CLK(clknet_4_2_0_clk),
    .D(\u_delay_line.dl_25 ),
    .RESET_B(net5),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\u_delay_line.data_24 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_24.u_inv_0  (.A(\u_delay_line.dl_24 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_24.dl_0 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_24.u_inv_1  (.A(\u_delay_line.u_dl_24.dl_0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_24.dl_1 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_24.u_inv_10  (.A(\u_delay_line.u_dl_24.dl_9 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_24.dl_10 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_24.u_inv_11  (.A(\u_delay_line.u_dl_24.dl_10 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.dl_25 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_24.u_inv_2  (.A(\u_delay_line.u_dl_24.dl_1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_24.dl_2 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_24.u_inv_3  (.A(\u_delay_line.u_dl_24.dl_2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_24.dl_3 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_24.u_inv_4  (.A(\u_delay_line.u_dl_24.dl_3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_24.dl_4 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_24.u_inv_5  (.A(\u_delay_line.u_dl_24.dl_4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_24.dl_5 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_24.u_inv_6  (.A(\u_delay_line.u_dl_24.dl_5 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_24.dl_6 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_24.u_inv_7  (.A(\u_delay_line.u_dl_24.dl_6 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_24.dl_7 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_24.u_inv_8  (.A(\u_delay_line.u_dl_24.dl_7 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_24.dl_8 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_24.u_inv_9  (.A(\u_delay_line.u_dl_24.dl_8 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_24.dl_9 ));
 sky130_fd_sc_hd__dfrtp_1 \u_delay_line.u_dl_25.u_ff  (.CLK(clknet_4_2_0_clk),
    .D(\u_delay_line.dl_26 ),
    .RESET_B(net5),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\u_delay_line.data_25 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_25.u_inv_0  (.A(\u_delay_line.dl_25 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_25.dl_0 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_25.u_inv_1  (.A(\u_delay_line.u_dl_25.dl_0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_25.dl_1 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_25.u_inv_10  (.A(\u_delay_line.u_dl_25.dl_9 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_25.dl_10 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_25.u_inv_11  (.A(\u_delay_line.u_dl_25.dl_10 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.dl_26 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_25.u_inv_2  (.A(\u_delay_line.u_dl_25.dl_1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_25.dl_2 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_25.u_inv_3  (.A(\u_delay_line.u_dl_25.dl_2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_25.dl_3 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_25.u_inv_4  (.A(\u_delay_line.u_dl_25.dl_3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_25.dl_4 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_25.u_inv_5  (.A(\u_delay_line.u_dl_25.dl_4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_25.dl_5 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_25.u_inv_6  (.A(\u_delay_line.u_dl_25.dl_5 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_25.dl_6 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_25.u_inv_7  (.A(\u_delay_line.u_dl_25.dl_6 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_25.dl_7 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_25.u_inv_8  (.A(\u_delay_line.u_dl_25.dl_7 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_25.dl_8 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_25.u_inv_9  (.A(\u_delay_line.u_dl_25.dl_8 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_25.dl_9 ));
 sky130_fd_sc_hd__dfrtp_1 \u_delay_line.u_dl_26.u_ff  (.CLK(clknet_4_2_0_clk),
    .D(\u_delay_line.dl_27 ),
    .RESET_B(net5),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\u_delay_line.data_26 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_26.u_inv_0  (.A(\u_delay_line.dl_26 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_26.dl_0 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_26.u_inv_1  (.A(\u_delay_line.u_dl_26.dl_0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_26.dl_1 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_26.u_inv_10  (.A(\u_delay_line.u_dl_26.dl_9 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_26.dl_10 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_26.u_inv_11  (.A(\u_delay_line.u_dl_26.dl_10 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.dl_27 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_26.u_inv_2  (.A(\u_delay_line.u_dl_26.dl_1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_26.dl_2 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_26.u_inv_3  (.A(\u_delay_line.u_dl_26.dl_2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_26.dl_3 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_26.u_inv_4  (.A(\u_delay_line.u_dl_26.dl_3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_26.dl_4 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_26.u_inv_5  (.A(\u_delay_line.u_dl_26.dl_4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_26.dl_5 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_26.u_inv_6  (.A(\u_delay_line.u_dl_26.dl_5 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_26.dl_6 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_26.u_inv_7  (.A(\u_delay_line.u_dl_26.dl_6 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_26.dl_7 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_26.u_inv_8  (.A(\u_delay_line.u_dl_26.dl_7 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_26.dl_8 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_26.u_inv_9  (.A(\u_delay_line.u_dl_26.dl_8 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_26.dl_9 ));
 sky130_fd_sc_hd__dfrtp_1 \u_delay_line.u_dl_27.u_ff  (.CLK(clknet_4_8_0_clk),
    .D(\u_delay_line.dl_28 ),
    .RESET_B(net11),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\u_delay_line.data_27 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_27.u_inv_0  (.A(\u_delay_line.dl_27 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_27.dl_0 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_27.u_inv_1  (.A(\u_delay_line.u_dl_27.dl_0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_27.dl_1 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_27.u_inv_10  (.A(\u_delay_line.u_dl_27.dl_9 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_27.dl_10 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_27.u_inv_11  (.A(\u_delay_line.u_dl_27.dl_10 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.dl_28 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_27.u_inv_2  (.A(\u_delay_line.u_dl_27.dl_1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_27.dl_2 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_27.u_inv_3  (.A(\u_delay_line.u_dl_27.dl_2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_27.dl_3 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_27.u_inv_4  (.A(\u_delay_line.u_dl_27.dl_3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_27.dl_4 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_27.u_inv_5  (.A(\u_delay_line.u_dl_27.dl_4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_27.dl_5 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_27.u_inv_6  (.A(\u_delay_line.u_dl_27.dl_5 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_27.dl_6 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_27.u_inv_7  (.A(\u_delay_line.u_dl_27.dl_6 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_27.dl_7 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_27.u_inv_8  (.A(\u_delay_line.u_dl_27.dl_7 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_27.dl_8 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_27.u_inv_9  (.A(\u_delay_line.u_dl_27.dl_8 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_27.dl_9 ));
 sky130_fd_sc_hd__dfrtp_1 \u_delay_line.u_dl_28.u_ff  (.CLK(clknet_4_8_0_clk),
    .D(\u_delay_line.dl_29 ),
    .RESET_B(net11),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\u_delay_line.data_28 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_28.u_inv_0  (.A(\u_delay_line.dl_28 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_28.dl_0 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_28.u_inv_1  (.A(\u_delay_line.u_dl_28.dl_0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_28.dl_1 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_28.u_inv_10  (.A(\u_delay_line.u_dl_28.dl_9 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_28.dl_10 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_28.u_inv_11  (.A(\u_delay_line.u_dl_28.dl_10 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.dl_29 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_28.u_inv_2  (.A(\u_delay_line.u_dl_28.dl_1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_28.dl_2 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_28.u_inv_3  (.A(\u_delay_line.u_dl_28.dl_2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_28.dl_3 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_28.u_inv_4  (.A(\u_delay_line.u_dl_28.dl_3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_28.dl_4 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_28.u_inv_5  (.A(\u_delay_line.u_dl_28.dl_4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_28.dl_5 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_28.u_inv_6  (.A(\u_delay_line.u_dl_28.dl_5 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_28.dl_6 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_28.u_inv_7  (.A(\u_delay_line.u_dl_28.dl_6 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_28.dl_7 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_28.u_inv_8  (.A(\u_delay_line.u_dl_28.dl_7 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_28.dl_8 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_28.u_inv_9  (.A(\u_delay_line.u_dl_28.dl_8 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_28.dl_9 ));
 sky130_fd_sc_hd__dfrtp_1 \u_delay_line.u_dl_29.u_ff  (.CLK(clknet_4_8_0_clk),
    .D(\u_delay_line.dl_30 ),
    .RESET_B(net11),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\u_delay_line.data_29 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_29.u_inv_0  (.A(\u_delay_line.dl_29 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_29.dl_0 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_29.u_inv_1  (.A(\u_delay_line.u_dl_29.dl_0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_29.dl_1 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_29.u_inv_10  (.A(\u_delay_line.u_dl_29.dl_9 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_29.dl_10 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_29.u_inv_11  (.A(\u_delay_line.u_dl_29.dl_10 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.dl_30 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_29.u_inv_2  (.A(\u_delay_line.u_dl_29.dl_1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_29.dl_2 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_29.u_inv_3  (.A(\u_delay_line.u_dl_29.dl_2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_29.dl_3 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_29.u_inv_4  (.A(\u_delay_line.u_dl_29.dl_3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_29.dl_4 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_29.u_inv_5  (.A(\u_delay_line.u_dl_29.dl_4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_29.dl_5 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_29.u_inv_6  (.A(\u_delay_line.u_dl_29.dl_5 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_29.dl_6 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_29.u_inv_7  (.A(\u_delay_line.u_dl_29.dl_6 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_29.dl_7 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_29.u_inv_8  (.A(\u_delay_line.u_dl_29.dl_7 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_29.dl_8 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_29.u_inv_9  (.A(\u_delay_line.u_dl_29.dl_8 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_29.dl_9 ));
 sky130_fd_sc_hd__dfrtp_2 \u_delay_line.u_dl_3.u_ff  (.CLK(clknet_4_0_0_clk),
    .D(\u_delay_line.dl_4 ),
    .RESET_B(net3),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\u_delay_line.data_3 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_3.u_inv_0  (.A(\u_delay_line.dl_3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_3.dl_0 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_3.u_inv_1  (.A(\u_delay_line.u_dl_3.dl_0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_3.dl_1 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_3.u_inv_10  (.A(\u_delay_line.u_dl_3.dl_9 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_3.dl_10 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_3.u_inv_11  (.A(\u_delay_line.u_dl_3.dl_10 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.dl_4 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_3.u_inv_2  (.A(\u_delay_line.u_dl_3.dl_1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_3.dl_2 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_3.u_inv_3  (.A(\u_delay_line.u_dl_3.dl_2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_3.dl_3 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_3.u_inv_4  (.A(\u_delay_line.u_dl_3.dl_3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_3.dl_4 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_3.u_inv_5  (.A(\u_delay_line.u_dl_3.dl_4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_3.dl_5 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_3.u_inv_6  (.A(\u_delay_line.u_dl_3.dl_5 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_3.dl_6 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_3.u_inv_7  (.A(\u_delay_line.u_dl_3.dl_6 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_3.dl_7 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_3.u_inv_8  (.A(\u_delay_line.u_dl_3.dl_7 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_3.dl_8 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_3.u_inv_9  (.A(\u_delay_line.u_dl_3.dl_8 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_3.dl_9 ));
 sky130_fd_sc_hd__dfrtp_1 \u_delay_line.u_dl_30.u_ff  (.CLK(clknet_4_10_0_clk),
    .D(\u_delay_line.dl_31 ),
    .RESET_B(net12),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\u_delay_line.data_30 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_30.u_inv_0  (.A(\u_delay_line.dl_30 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_30.dl_0 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_30.u_inv_1  (.A(\u_delay_line.u_dl_30.dl_0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_30.dl_1 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_30.u_inv_10  (.A(\u_delay_line.u_dl_30.dl_9 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_30.dl_10 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_30.u_inv_11  (.A(\u_delay_line.u_dl_30.dl_10 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.dl_31 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_30.u_inv_2  (.A(\u_delay_line.u_dl_30.dl_1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_30.dl_2 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_30.u_inv_3  (.A(\u_delay_line.u_dl_30.dl_2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_30.dl_3 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_30.u_inv_4  (.A(\u_delay_line.u_dl_30.dl_3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_30.dl_4 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_30.u_inv_5  (.A(\u_delay_line.u_dl_30.dl_4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_30.dl_5 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_30.u_inv_6  (.A(\u_delay_line.u_dl_30.dl_5 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_30.dl_6 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_30.u_inv_7  (.A(\u_delay_line.u_dl_30.dl_6 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_30.dl_7 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_30.u_inv_8  (.A(\u_delay_line.u_dl_30.dl_7 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_30.dl_8 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_30.u_inv_9  (.A(\u_delay_line.u_dl_30.dl_8 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_30.dl_9 ));
 sky130_fd_sc_hd__dfrtp_1 \u_delay_line.u_dl_31.u_ff  (.CLK(clknet_4_8_0_clk),
    .D(\u_delay_line.dl_32 ),
    .RESET_B(net11),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\u_delay_line.data_31 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_31.u_inv_0  (.A(\u_delay_line.dl_31 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_31.dl_0 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_31.u_inv_1  (.A(\u_delay_line.u_dl_31.dl_0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_31.dl_1 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_31.u_inv_10  (.A(\u_delay_line.u_dl_31.dl_9 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_31.dl_10 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_31.u_inv_11  (.A(\u_delay_line.u_dl_31.dl_10 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.dl_32 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_31.u_inv_2  (.A(\u_delay_line.u_dl_31.dl_1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_31.dl_2 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_31.u_inv_3  (.A(\u_delay_line.u_dl_31.dl_2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_31.dl_3 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_31.u_inv_4  (.A(\u_delay_line.u_dl_31.dl_3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_31.dl_4 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_31.u_inv_5  (.A(\u_delay_line.u_dl_31.dl_4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_31.dl_5 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_31.u_inv_6  (.A(\u_delay_line.u_dl_31.dl_5 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_31.dl_6 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_31.u_inv_7  (.A(\u_delay_line.u_dl_31.dl_6 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_31.dl_7 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_31.u_inv_8  (.A(\u_delay_line.u_dl_31.dl_7 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_31.dl_8 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_31.u_inv_9  (.A(\u_delay_line.u_dl_31.dl_8 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_31.dl_9 ));
 sky130_fd_sc_hd__dfrtp_1 \u_delay_line.u_dl_4.u_ff  (.CLK(clknet_4_0_0_clk),
    .D(\u_delay_line.dl_5 ),
    .RESET_B(net3),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\u_delay_line.data_4 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_4.u_inv_0  (.A(\u_delay_line.dl_4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_4.dl_0 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_4.u_inv_1  (.A(\u_delay_line.u_dl_4.dl_0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_4.dl_1 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_4.u_inv_10  (.A(\u_delay_line.u_dl_4.dl_9 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_4.dl_10 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_4.u_inv_11  (.A(\u_delay_line.u_dl_4.dl_10 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.dl_5 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_4.u_inv_2  (.A(\u_delay_line.u_dl_4.dl_1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_4.dl_2 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_4.u_inv_3  (.A(\u_delay_line.u_dl_4.dl_2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_4.dl_3 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_4.u_inv_4  (.A(\u_delay_line.u_dl_4.dl_3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_4.dl_4 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_4.u_inv_5  (.A(\u_delay_line.u_dl_4.dl_4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_4.dl_5 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_4.u_inv_6  (.A(\u_delay_line.u_dl_4.dl_5 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_4.dl_6 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_4.u_inv_7  (.A(\u_delay_line.u_dl_4.dl_6 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_4.dl_7 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_4.u_inv_8  (.A(\u_delay_line.u_dl_4.dl_7 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_4.dl_8 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_4.u_inv_9  (.A(\u_delay_line.u_dl_4.dl_8 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_4.dl_9 ));
 sky130_fd_sc_hd__dfrtp_2 \u_delay_line.u_dl_5.u_ff  (.CLK(clknet_4_0_0_clk),
    .D(\u_delay_line.dl_6 ),
    .RESET_B(net4),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\u_delay_line.data_5 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_5.u_inv_0  (.A(\u_delay_line.dl_5 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_5.dl_0 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_5.u_inv_1  (.A(\u_delay_line.u_dl_5.dl_0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_5.dl_1 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_5.u_inv_10  (.A(\u_delay_line.u_dl_5.dl_9 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_5.dl_10 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_5.u_inv_11  (.A(\u_delay_line.u_dl_5.dl_10 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.dl_6 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_5.u_inv_2  (.A(\u_delay_line.u_dl_5.dl_1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_5.dl_2 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_5.u_inv_3  (.A(\u_delay_line.u_dl_5.dl_2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_5.dl_3 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_5.u_inv_4  (.A(\u_delay_line.u_dl_5.dl_3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_5.dl_4 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_5.u_inv_5  (.A(\u_delay_line.u_dl_5.dl_4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_5.dl_5 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_5.u_inv_6  (.A(\u_delay_line.u_dl_5.dl_5 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_5.dl_6 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_5.u_inv_7  (.A(\u_delay_line.u_dl_5.dl_6 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_5.dl_7 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_5.u_inv_8  (.A(\u_delay_line.u_dl_5.dl_7 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_5.dl_8 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_5.u_inv_9  (.A(\u_delay_line.u_dl_5.dl_8 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_5.dl_9 ));
 sky130_fd_sc_hd__dfrtp_1 \u_delay_line.u_dl_6.u_ff  (.CLK(clknet_4_1_0_clk),
    .D(\u_delay_line.dl_7 ),
    .RESET_B(net4),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\u_delay_line.data_6 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_6.u_inv_0  (.A(\u_delay_line.dl_6 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_6.dl_0 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_6.u_inv_1  (.A(\u_delay_line.u_dl_6.dl_0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_6.dl_1 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_6.u_inv_10  (.A(\u_delay_line.u_dl_6.dl_9 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_6.dl_10 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_6.u_inv_11  (.A(\u_delay_line.u_dl_6.dl_10 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.dl_7 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_6.u_inv_2  (.A(\u_delay_line.u_dl_6.dl_1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_6.dl_2 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_6.u_inv_3  (.A(\u_delay_line.u_dl_6.dl_2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_6.dl_3 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_6.u_inv_4  (.A(\u_delay_line.u_dl_6.dl_3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_6.dl_4 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_6.u_inv_5  (.A(\u_delay_line.u_dl_6.dl_4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_6.dl_5 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_6.u_inv_6  (.A(\u_delay_line.u_dl_6.dl_5 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_6.dl_6 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_6.u_inv_7  (.A(\u_delay_line.u_dl_6.dl_6 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_6.dl_7 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_6.u_inv_8  (.A(\u_delay_line.u_dl_6.dl_7 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_6.dl_8 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_6.u_inv_9  (.A(\u_delay_line.u_dl_6.dl_8 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_6.dl_9 ));
 sky130_fd_sc_hd__dfrtp_2 \u_delay_line.u_dl_7.u_ff  (.CLK(clknet_4_4_0_clk),
    .D(\u_delay_line.dl_8 ),
    .RESET_B(net7),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\u_delay_line.data_7 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_7.u_inv_0  (.A(\u_delay_line.dl_7 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_7.dl_0 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_7.u_inv_1  (.A(\u_delay_line.u_dl_7.dl_0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_7.dl_1 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_7.u_inv_10  (.A(\u_delay_line.u_dl_7.dl_9 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_7.dl_10 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_7.u_inv_11  (.A(\u_delay_line.u_dl_7.dl_10 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.dl_8 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_7.u_inv_2  (.A(\u_delay_line.u_dl_7.dl_1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_7.dl_2 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_7.u_inv_3  (.A(\u_delay_line.u_dl_7.dl_2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_7.dl_3 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_7.u_inv_4  (.A(\u_delay_line.u_dl_7.dl_3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_7.dl_4 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_7.u_inv_5  (.A(\u_delay_line.u_dl_7.dl_4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_7.dl_5 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_7.u_inv_6  (.A(\u_delay_line.u_dl_7.dl_5 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_7.dl_6 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_7.u_inv_7  (.A(\u_delay_line.u_dl_7.dl_6 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_7.dl_7 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_7.u_inv_8  (.A(\u_delay_line.u_dl_7.dl_7 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_7.dl_8 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_7.u_inv_9  (.A(\u_delay_line.u_dl_7.dl_8 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_7.dl_9 ));
 sky130_fd_sc_hd__dfrtp_1 \u_delay_line.u_dl_8.u_ff  (.CLK(clknet_4_4_0_clk),
    .D(\u_delay_line.dl_9 ),
    .RESET_B(net7),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\u_delay_line.data_8 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_8.u_inv_0  (.A(\u_delay_line.dl_8 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_8.dl_0 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_8.u_inv_1  (.A(\u_delay_line.u_dl_8.dl_0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_8.dl_1 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_8.u_inv_10  (.A(\u_delay_line.u_dl_8.dl_9 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_8.dl_10 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_8.u_inv_11  (.A(\u_delay_line.u_dl_8.dl_10 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.dl_9 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_8.u_inv_2  (.A(\u_delay_line.u_dl_8.dl_1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_8.dl_2 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_8.u_inv_3  (.A(\u_delay_line.u_dl_8.dl_2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_8.dl_3 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_8.u_inv_4  (.A(\u_delay_line.u_dl_8.dl_3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_8.dl_4 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_8.u_inv_5  (.A(\u_delay_line.u_dl_8.dl_4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_8.dl_5 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_8.u_inv_6  (.A(\u_delay_line.u_dl_8.dl_5 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_8.dl_6 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_8.u_inv_7  (.A(\u_delay_line.u_dl_8.dl_6 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_8.dl_7 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_8.u_inv_8  (.A(\u_delay_line.u_dl_8.dl_7 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_8.dl_8 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_8.u_inv_9  (.A(\u_delay_line.u_dl_8.dl_8 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_8.dl_9 ));
 sky130_fd_sc_hd__dfrtp_1 \u_delay_line.u_dl_9.u_ff  (.CLK(clknet_4_4_0_clk),
    .D(\u_delay_line.dl_10 ),
    .RESET_B(net7),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\u_delay_line.data_9 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_9.u_inv_0  (.A(\u_delay_line.dl_9 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_9.dl_0 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_9.u_inv_1  (.A(\u_delay_line.u_dl_9.dl_0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_9.dl_1 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_9.u_inv_10  (.A(\u_delay_line.u_dl_9.dl_9 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_9.dl_10 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_9.u_inv_11  (.A(\u_delay_line.u_dl_9.dl_10 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.dl_10 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_9.u_inv_2  (.A(\u_delay_line.u_dl_9.dl_1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_9.dl_2 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_9.u_inv_3  (.A(\u_delay_line.u_dl_9.dl_2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_9.dl_3 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_9.u_inv_4  (.A(\u_delay_line.u_dl_9.dl_3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_9.dl_4 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_9.u_inv_5  (.A(\u_delay_line.u_dl_9.dl_4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_9.dl_5 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_9.u_inv_6  (.A(\u_delay_line.u_dl_9.dl_5 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_9.dl_6 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_9.u_inv_7  (.A(\u_delay_line.u_dl_9.dl_6 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_9.dl_7 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_9.u_inv_8  (.A(\u_delay_line.u_dl_9.dl_7 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_9.dl_8 ));
 sky130_fd_sc_hd__inv_2 \u_delay_line.u_dl_9.u_inv_9  (.A(\u_delay_line.u_dl_9.dl_8 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_delay_line.u_dl_9.dl_9 ));
 sky130_fd_sc_hd__inv_1 \u_delay_line.u_inv_0  (.A(\u_delay_line.dl_32 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 assign uio_oe[0] = net20;
 assign uio_oe[1] = net21;
 assign uio_oe[2] = net22;
 assign uio_oe[3] = net23;
 assign uio_oe[4] = net24;
 assign uio_oe[5] = net25;
 assign uio_oe[6] = net26;
 assign uio_oe[7] = net27;
 assign uio_out[0] = net28;
 assign uio_out[1] = net29;
 assign uio_out[2] = net30;
 assign uio_out[3] = net31;
 assign uio_out[4] = net32;
 assign uio_out[5] = net33;
 assign uio_out[6] = net34;
 assign uio_out[7] = net35;
 assign uo_out[1] = net36;
 assign uo_out[2] = net37;
 assign uo_out[3] = net38;
 assign uo_out[4] = net39;
 assign uo_out[5] = net40;
 assign uo_out[6] = net41;
 assign uo_out[7] = net42;
endmodule
